`define PHY_PORT_TABLE_CONTENT         reg_config.phy_port_table.table_index
`define LOGIC_PORT_TABLE_CONTENT       reg_config.logic_port_table.table_index
`define L2_PROTOCOL_TABLE_CONTENT      reg_config.l2_protocol_table.table_index
`define IPHB_TABLE_CONTENT             reg_config.iphb_table.table_index
`define IVLAN_XLATE_TABLE_CONTENT      reg_config.ivlan_xlate_table.table_index
`define IVLAN_PROPERTY_TABLE_CONTENT   reg_config.ivlan_property_table.table_index
`define IVLAN_ACTION_TABLE_CONTENT     reg_config.ivlan_action_table.table_index
`define IVLAN_STG_TABLE_CONTENT        reg_config.ivlan_stg_table.table_index
`define L2_MAC_TABLE_CONTENT           reg_config.l2_mac_table.table_index
`define STORM_POLICER_ID_TABLE_CONTENT reg_config.storm_policer_id_table.table_index
`define ING_FLOW_TABLE_CONTENT         reg_config.ing_flow_table.table_index
`define ING_FLOW_PRO_TABLE_CONTENT     reg_config.ing_flow_pro_table.table_index
`define ING_GATE_TABLE_CONTENT         reg_config.ing_gate_table.table_index
`define POLICER_CONF_TABLE_CONTENT     reg_config.policer_conf_table.table_index
`define POLICER_TOKEN_TABLE_CONTENT    reg_config.policer_token_table.table_index
`define FRER_REC_TABLE_CONTENT         reg_config.frer_rec_table.table_index
`define RX_PTP_FORWARD_TABLE_CONTENT   reg_config.rx_ptp_forward_table.table_index
`define OUT_FP_TABLE_CONTENT           reg_config.out_fp_table.table_index
`define L2_MC_TABLE_CONTENT            reg_config.l2_mc_table.table_index
`define TIME_SLOT_TABLE_CONTENT        reg_config.time_slot_table.table_index
`define EVLAN_XLATE_TABLE_CONTENT      reg_config.evlan_xlate_table.table_index
`define EVLAN_ACTION_TABLE_CONTENT     reg_config.evlan_action_table.table_index
`define EVLAN_PROPERTY_TABLE_CONTENT   reg_config.evlan_property_table.table_index
`define EVLAN_STG_TABLE_CONTENT        reg_config.evlan_stg_table.table_index
`define OPORT_PRO_TABLE_CONTENT        reg_config.oport_pro_table.table_index
`define DOT1P_MAP_TABLE_CONTENT        reg_config.dot1p_map_table.table_index
`define LAG_SEL_PORT_TABLE_CONTENT     reg_config.lag_sel_port_table.table_index
`define O_PHY_PORT_PRO_TABLE_CONTENT   reg_config.o_phy_port_pro_table.table_index
`define GATHER_INIT_TABLE_CONTENT      reg_config.gather_init_table.table_index

`define BASE_OFFSET   15'b100_0000_0000_0000
`define BASE_OFFSET_GATHER   16'b011_0000_0000_0000
`define PP_VER_YEAR	        (`BASE_OFFSET+'h0000)
`define PP_VER_MONTH_DAY	(`BASE_OFFSET+'h0002)
`define PP_VER_HOUR_MIN	    (`BASE_OFFSET+'h0004)
`define PP_TEST_REG	        (`BASE_OFFSET+'h0006)	
// PHY_PORT_TABLE	
`define PHY_PORT_TABLE_STATUS	(`BASE_OFFSET+'h0020)	
`define PHY_PORT_TABLE_CONTROL	(`BASE_OFFSET+'h0022)	
`define PHY_PORT_TABLE_DIN_0	(`BASE_OFFSET+'h0024)	
`define PHY_PORT_TABLE_DIN_1	(`BASE_OFFSET+'h0026)
`define PHY_PORT_TABLE_DIN_2	(`BASE_OFFSET+'h0028)
`define PHY_PORT_TABLE_DIN_3	(`BASE_OFFSET+'h002A)
`define PHY_PORT_TABLE_DIN_4	(`BASE_OFFSET+'h002C)
`define PHY_PORT_TABLE_DIN_5	(`BASE_OFFSET+'h002E)
`define PHY_PORT_TABLE_DIN_6	(`BASE_OFFSET+'h0030)
`define PHY_PORT_TABLE_DOUT_0	(`BASE_OFFSET+'h0032)	
`define PHY_PORT_TABLE_DOUT_1	(`BASE_OFFSET+'h0034)
`define PHY_PORT_TABLE_DOUT_2	(`BASE_OFFSET+'h0036)
`define PHY_PORT_TABLE_DOUT_3	(`BASE_OFFSET+'h0038)
`define PHY_PORT_TABLE_DOUT_4	(`BASE_OFFSET+'h003A)
`define PHY_PORT_TABLE_DOUT_5	(`BASE_OFFSET+'h003C)
`define PHY_PORT_TABLE_DOUT_6	(`BASE_OFFSET+'h003E)	
// LOGIC_PORT_TABLE	
`define LOGIC_PORT_TABLE_STATUS	 (`BASE_OFFSET+'h0200)	
`define LOGIC_PORT_TABLE_CONTROL (`BASE_OFFSET+'h0202)	
`define LOGIC_PORT_TABLE_DIN_0	 (`BASE_OFFSET+'h0204)	
`define LOGIC_PORT_TABLE_DIN_1	 (`BASE_OFFSET+'h0206)
`define LOGIC_PORT_TABLE_DIN_2	 (`BASE_OFFSET+'h0208)
`define LOGIC_PORT_TABLE_DIN_3	 (`BASE_OFFSET+'h020A)
`define LOGIC_PORT_TABLE_DIN_4	 (`BASE_OFFSET+'h020C)
`define LOGIC_PORT_TABLE_DIN_5	 (`BASE_OFFSET+'h020E)
`define LOGIC_PORT_TABLE_DIN_6	 (`BASE_OFFSET+'h0210)
`define LOGIC_PORT_TABLE_DIN_7	 (`BASE_OFFSET+'h0212)
`define LOGIC_PORT_TABLE_DOUT_0	 (`BASE_OFFSET+'h0214)	
`define LOGIC_PORT_TABLE_DOUT_1	 (`BASE_OFFSET+'h0216)
`define LOGIC_PORT_TABLE_DOUT_2	 (`BASE_OFFSET+'h0218)
`define LOGIC_PORT_TABLE_DOUT_3	 (`BASE_OFFSET+'h021A)
`define LOGIC_PORT_TABLE_DOUT_4	 (`BASE_OFFSET+'h021C)
`define LOGIC_PORT_TABLE_DOUT_5	 (`BASE_OFFSET+'h021E)
`define LOGIC_PORT_TABLE_DOUT_6	 (`BASE_OFFSET+'h0220)
`define LOGIC_PORT_TABLE_DOUT_7	 (`BASE_OFFSET+'h0222)
// L2_PROTOCOL_TABLE	
`define L2_PROTOCOL_TABLE_STATUS	(`BASE_OFFSET+'h0240)	
`define L2_PROTOCOL_TABLE_CONTROL	(`BASE_OFFSET+'h0242)	
`define L2_PROTOCOL_TABLE_DIN_0	    (`BASE_OFFSET+'h0244)	
`define L2_PROTOCOL_TABLE_DIN_1	    (`BASE_OFFSET+'h0246)
`define L2_PROTOCOL_TABLE_DOUT_0	(`BASE_OFFSET+'h0248)	
`define L2_PROTOCOL_TABLE_DOUT_1	(`BASE_OFFSET+'h024a)	
`define PAUSE_PCKT_DROP_EN	        (`BASE_OFFSET+'h0400)	
`define CRC_ERR_DROP_R_TRIG	        (`BASE_OFFSET+'h0402)	
`define CRC_ERR_DROP_ROUT_H	        (`BASE_OFFSET+'h0404)	
`define CRC_ERR_DROP_ROUT_L	        (`BASE_OFFSET+'h0406)
`define BIND_SA_DROP_R_TRIG	        (`BASE_OFFSET+'h0408)	
`define BIND_SA_DROP_ROUT_H	        (`BASE_OFFSET+'h040A)	
`define BIND_SA_DROP_ROUT_L	        (`BASE_OFFSET+'h040C)
`define L2_CTL_DROP_R_TRIG	        (`BASE_OFFSET+'h040E)	
`define L2_CTL_DROP_ROUT_H	        (`BASE_OFFSET+'h0410)	
`define L2_CTL_DROP_ROUT_L	        (`BASE_OFFSET+'h0412)
`define TPID_REG_0	                (`BASE_OFFSET+'h0420)
`define TPID_REG_1	                (`BASE_OFFSET+'h0422)
`define TPID_REG_2	                (`BASE_OFFSET+'h0424)
`define TPID_REG_3	                (`BASE_OFFSET+'h0426)	
// IPHB_TABLE	
`define IPHB_TABLE_STATUS	(`BASE_OFFSET+'h0600)	
`define IPHB_TABLE_CONTROL	(`BASE_OFFSET+'h0602)
`define IPHB_T_CONF_DIN	    (`BASE_OFFSET+'h0604)	
`define IPHB_T_CONF_DOUT	(`BASE_OFFSET+'h0606)	
// IVLAN_XLATE_TABLE	
`define IVLAN_XLATE_TABLE_STATUS	(`BASE_OFFSET+'h060A)	
`define IVLAN_XLATE_TABLE_CONTROL	(`BASE_OFFSET+'h060C)
`define IVLAN_XLATE_T_CONF_KEY	    (`BASE_OFFSET+'h060E)
`define IVLAN_XLATE_T_CONF_DIN_0	(`BASE_OFFSET+'h0610)	
`define IVLAN_XLATE_T_CONF_DIN_1	(`BASE_OFFSET+'h0612)
`define IVLAN_XLATE_T_CONF_DOUT_0	(`BASE_OFFSET+'h0614)
`define IVLAN_XLATE_T_CONF_DOUT_1	(`BASE_OFFSET+'h0616)
`define IVLAN_XLATE_T_CONF_DOUT_2	(`BASE_OFFSET+'h0618)
// IVLAN_PROPERTY_TABLE	
`define IVLAN_PROPERTY_TABLE_STATUS	    (`BASE_OFFSET+'h0620)	
`define IVLAN_PROPERTY_TABLE_CONTROL	(`BASE_OFFSET+'h0622)
`define IVLAN_PROPERTY_T_CONF_DIN_0	    (`BASE_OFFSET+'h0624)
`define IVLAN_PROPERTY_T_CONF_DIN_1	    (`BASE_OFFSET+'h0626)
`define IVLAN_PROPERTY_T_CONF_DIN_2	    (`BASE_OFFSET+'h0628)
`define IVLAN_PROPERTY_T_CONF_DIN_3	    (`BASE_OFFSET+'h062A)
`define IVLAN_PROPERTY_T_CONF_DOUT_0	(`BASE_OFFSET+'h062C)
`define IVLAN_PROPERTY_T_CONF_DOUT_1	(`BASE_OFFSET+'h062E)
`define IVLAN_PROPERTY_T_CONF_DOUT_2	(`BASE_OFFSET+'h0630)
`define IVLAN_PROPERTY_T_CONF_DOUT_3	(`BASE_OFFSET+'h0632)
// IVLAN_ACTION_TABLE	
`define IVLAN_ACTION_TABLE_STATUS	(`BASE_OFFSET+'h0640)	
`define IVLAN_ACTION_TABLE_CONTROL	(`BASE_OFFSET+'h0642)
`define IVLAN_ACTION_T_CONF_DIN_0	(`BASE_OFFSET+'h0644)
`define IVLAN_ACTION_T_CONF_DIN_1	(`BASE_OFFSET+'h0646)
`define IVLAN_ACTION_T_CONF_DOUT_0	(`BASE_OFFSET+'h0648)
`define IVLAN_ACTION_T_CONF_DOUT_1	(`BASE_OFFSET+'h064A)
// IVLAN_STG_TABLE	
`define IVLAN_STG_TABLE_STATUS	(`BASE_OFFSET+'h0660)	
`define IVLAN_STG_TABLE_CONTROL	(`BASE_OFFSET+'h0662)	
`define ISTG_T_CONF_DIN_0	    (`BASE_OFFSET+'h0664)
`define ISTG_T_CONF_DIN_1	    (`BASE_OFFSET+'h0666)
`define ISTG_T_CONF_DIN_2	    (`BASE_OFFSET+'h0668)
`define ISTG_T_CONF_DIN_3	    (`BASE_OFFSET+'h066A)
`define ISTG_T_CONF_DOUT_0	    (`BASE_OFFSET+'h066C)
`define ISTG_T_CONF_DOUT_1	    (`BASE_OFFSET+'h066E)
`define ISTG_T_CONF_DOUT_2	    (`BASE_OFFSET+'h0670)
`define ISTG_T_CONF_DOUT_3	    (`BASE_OFFSET+'h0672)
`define VT_MISS_DROP_R_TRIG	    (`BASE_OFFSET+'h0680)
`define VT_MISS_DROP_ROUT_H	    (`BASE_OFFSET+'h0682)	
`define VT_MISS_DROP_ROUT_L	    (`BASE_OFFSET+'h0684)
`define VLAN_FILTER_DROP_R_TRIG	(`BASE_OFFSET+'h0686)	
`define VLAN_FILTER_DROP_ROUT_H	(`BASE_OFFSET+'h0688)
`define VLAN_FILTER_DROP_ROUT_1	(`BASE_OFFSET+'h068A)
`define STP_DROP_R_TRIG	        (`BASE_OFFSET+'h068C)
`define STP_DROP_ROUT_H	        (`BASE_OFFSET+'h068E)
`define STP_DROP_ROUT_L	        (`BASE_OFFSET+'h0690)
// L2_MAC_TABLE	
`define L2_MAC_TABLE_STATUS	    (`BASE_OFFSET+'h0800)
`define L2_MAC_TABLE_CONTROL	(`BASE_OFFSET+'h0802)
`define L2M_T_CONF_KEY_0	    (`BASE_OFFSET+'h0804)
`define L2M_T_CONF_KEY_1	    (`BASE_OFFSET+'h0806)
`define L2M_T_CONF_KEY_2	    (`BASE_OFFSET+'h0808)
`define L2M_T_CONF_DIN_0	    (`BASE_OFFSET+'h080A)	
`define L2M_T_CONF_DIN_1	    (`BASE_OFFSET+'h080C)
`define L2M_T_CONF_DOUT_0	    (`BASE_OFFSET+'h080E)
`define L2M_T_CONF_DOUT_1	    (`BASE_OFFSET+'h0810)
`define L2M_T_CONF_DOUT_2	    (`BASE_OFFSET+'h0812)
`define L2M_T_CONF_DOUT_3	    (`BASE_OFFSET+'h0814)
`define L2M_T_CONF_DOUT_4	    (`BASE_OFFSET+'h0816)
`define L2MT_AGE_TIMER_H	    (`BASE_OFFSET+'h0818)	
`define L2MT_AGE_TIMER_L	    (`BASE_OFFSET+'h081A)
`define IP_BIND_DROP_R_TRIG	    (`BASE_OFFSET+'h0820)	
`define IP_BIND_DROP_ROUT_H	    (`BASE_OFFSET+'h0822)	
`define IP_BIND_DROP_ROUT_L	    (`BASE_OFFSET+'h0824)	
`define L2_SRC_DROP_R_TRIG	    (`BASE_OFFSET+'h0826)	
`define L2_SRC_DROP_ROUT_H	    (`BASE_OFFSET+'h0828)	
`define L2_SRC_DROP_ROUT_L	    (`BASE_OFFSET+'h082A)	
`define L2_DST_DROP_R_TRIG	    (`BASE_OFFSET+'h082C)	
`define L2_DST_DROP_ROUT_H	    (`BASE_OFFSET+'h082E)
`define L2_DST_DROP_ROUT_L	    (`BASE_OFFSET+'h0830)
//`define STORM_POLICER_ID_TABLE	
`define STORM_POLICER_ID_TABLE_STATUS	(`BASE_OFFSET+'h0A00)	
`define STORM_POLICER_ID_TABLE_CONTROL	(`BASE_OFFSET+'h0A02)	
`define STORM_PID_T_CONF_DIN_0	        (`BASE_OFFSET+'h0A04)	
`define STORM_PID_T_CONF_DIN_1	        (`BASE_OFFSET+'h0A06)
`define STORM_PID_T_CONF_DOUT_0	        (`BASE_OFFSET+'h0A08)	
`define STORM_PID_T_CONF_DOUT_1	        (`BASE_OFFSET+'h0A0A)
//ING_FLOW_TABLE	
`define ING_FLOW_TABLE_STATUS	(`BASE_OFFSET+'h0A20)
`define ING_FLOW_TABLE_CONTROL	(`BASE_OFFSET+'h0A22)	
`define ING_FLOW_T_CONF_KEY_0	(`BASE_OFFSET+'h0A24)
`define ING_FLOW_T_CONF_KEY_1	(`BASE_OFFSET+'h0A26)
`define ING_FLOW_T_CONF_KEY_2	(`BASE_OFFSET+'h0A28)
`define ING_FLOW_T_CONF_KEY_3	(`BASE_OFFSET+'h0A2A)
`define ING_FLOW_T_CONF_DIN	    (`BASE_OFFSET+'h0A2C)	
`define ING_FLOW_T_CONF_DOUT_0	(`BASE_OFFSET+'h0A2E)
`define ING_FLOW_T_CONF_DOUT_1	(`BASE_OFFSET+'h0A30)
`define ING_FLOW_T_CONF_DOUT_2	(`BASE_OFFSET+'h0A32)
`define ING_FLOW_T_CONF_DOUT_3	(`BASE_OFFSET+'h0A34)
`define ING_FLOW_T_CONF_DOUT_4	(`BASE_OFFSET+'h0A36)
// ING_FLOW_PRO_TABLE	
`define ING_FLOW_PRO_TABLE_STATUS	(`BASE_OFFSET+'h0A40)	
`define ING_FLOW_PRO_TABLE_CONTROL	(`BASE_OFFSET+'h0A42)	
`define ING_FLOW_PRO_T_CONF_DIN_0	(`BASE_OFFSET+'h0A44)	
`define ING_FLOW_PRO_T_CONF_DIN_2	(`BASE_OFFSET+'h0A46)
`define ING_FLOW_PRO_T_CONF_DOUT_0	(`BASE_OFFSET+'h0A48)	
`define ING_FLOW_PRO_T_CONF_DOUT_1	(`BASE_OFFSET+'h0A4A)
// ING_GATE_TABLE	
`define ING_GATE_TABLE_STATUS	(`BASE_OFFSET+'h0A60)	
`define ING_GATE_TABLE_CONTROL	(`BASE_OFFSET+'h0A62)	
`define ING_GATE_T_CONF_DIN_0	(`BASE_OFFSET+'h0A64)	
`define ING_GATE_T_CONF_DIN_1	(`BASE_OFFSET+'h0A66)
`define ING_GATE_T_CONF_DOUT_0	(`BASE_OFFSET+'h0A68)	
`define ING_GATE_T_CONF_DOUT_1	(`BASE_OFFSET+'h0A6A)
//`define POLICER_CONF_TABLE	
`define POLICER_CONF_TABLE_STATUS	(`BASE_OFFSET+'h0A80)
`define POLICER_CONF_TABLE_CONTROL	(`BASE_OFFSET+'h0A82)	
`define POLICER_C_T_CONF_DIN_0	    (`BASE_OFFSET+'h0A84)	
`define POLICER_C_T_CONF_DIN_1	    (`BASE_OFFSET+'h0A86)
`define POLICER_C_T_CONF_DIN_2	    (`BASE_OFFSET+'h0A88)
`define POLICER_C_T_CONF_DOUT_0	    (`BASE_OFFSET+'h0A8A)	
`define POLICER_C_T_CONF_DOUT_1	    (`BASE_OFFSET+'h0A8C)
`define POLICER_C_T_CONF_DOUT_2	    (`BASE_OFFSET+'h0A8E)
`define POLICER_TIMER_REG	        (`BASE_OFFSET+'h0A90)
// POLICER_TOKEN_TABLE	
`define POLICER_TOKEN_TABLE_STATUS	(`BASE_OFFSET+'h0AA0)	
`define POLICER_TOKEN_TABLE_CONTROL	(`BASE_OFFSET+'h0AA2)
`define POLICER_TOKEN_T_CONF_DIN_0	(`BASE_OFFSET+'h0AA4)
`define POLICER_TOKEN_T_CONF_DIN_1	(`BASE_OFFSET+'h0AA6)
`define POLICER_TOKEN_T_CONF_DOUT_0	(`BASE_OFFSET+'h0AA8)
`define POLICER_TOKEN_T_CONF_DOUT_1	(`BASE_OFFSET+'h0AAA)
`define ING_GATE_DROP_R_TRIG	    (`BASE_OFFSET+'h0AC0)	
`define ING_GATE_DROP_ROUT_H	    (`BASE_OFFSET+'h0AC2)	
`define ING_GATE_DROP_ROUT_L	    (`BASE_OFFSET+'h0AC4)
`define ING_POLICER_DROP_R_TRIG	    (`BASE_OFFSET+'h0AC6)	
`define ING_POLICER_DROP_ROUT_H	    (`BASE_OFFSET+'h0AC8)	
`define ING_POLICER_DROP_ROUT_L	    (`BASE_OFFSET+'h0ACA)	
// TIME_SLOT_RAM	
`define TIME_SLOT_RAM_STATUS	(`BASE_OFFSET+'h0AE0)	
`define TIME_SLOT_RAM_CONTROL	(`BASE_OFFSET+'h0AE2)	
`define CONF_SLOT_RAM_WDATA_0	(`BASE_OFFSET+'h0AE4)
`define CONF_SLOT_RAM_WDATA_1	(`BASE_OFFSET+'h0AE6)
`define CONF_SLOT_RAM_RDATA_0	(`BASE_OFFSET+'h0AE8)
`define CONF_SLOT_RAM_RDATA_1	(`BASE_OFFSET+'h0AEA)
`define ADMIN_BASE_TIME_0	    (`BASE_OFFSET+'h0AEC)
`define ADMIN_BASE_TIME_1	    (`BASE_OFFSET+'h0AEE)
`define ADMIN_BASE_TIME_2	    (`BASE_OFFSET+'h0AF0)
`define ADMIN_BASE_TIME_3	    (`BASE_OFFSET+'h0AF2)	
`define ADMIN_CYCLE_TIME_0	    (`BASE_OFFSET+'h0AF4)
`define ADMIN_CYCLE_TIME_1	    (`BASE_OFFSET+'h0AF6)
`define ADMIN_CYCLE_TIME_2	    (`BASE_OFFSET+'h0AF8)
`define ADMIN_CYCLE_TIME_3	    (`BASE_OFFSET+'h0AFA)	
`define ADMIN_SLOT_NUM	                (`BASE_OFFSET+'h0AFC)	
`define TIME_SLOT_CONF_CONTROL_STATUS	(`BASE_OFFSET+'h0AFE)	
`define OPER_BASE_TIME_0	(`BASE_OFFSET+'h0B00)
`define OPER_BASE_TIME_1	(`BASE_OFFSET+'h0B02)
`define OPER_BASE_TIME_2	(`BASE_OFFSET+'h0B04)
`define OPER_BASE_TIME_3	(`BASE_OFFSET+'h0B06)
`define OPER_CYCLE_TIME_0	(`BASE_OFFSET+'h0B08)
`define OPER_CYCLE_TIME_1	(`BASE_OFFSET+'h0B0A)
`define OPER_CYCLE_TIME_2	(`BASE_OFFSET+'h0B0C)
`define OPER_CYCLE_TIME_3	(`BASE_OFFSET+'h0B0E)
`define OPER_SLOT_NUM	    (`BASE_OFFSET+'h0B10)
// FRER_REC_TABLE	
`define FRER_REC_TABLE_STATUS	(`BASE_OFFSET+'h0C00)	
`define FRER_REC_TABLE_CONTROL	(`BASE_OFFSET+'h0C02)	
`define FRER_REC_T_CONF_DIN_0	(`BASE_OFFSET+'h0C04)
`define FRER_REC_T_CONF_DIN_1	(`BASE_OFFSET+'h0C06)
`define FRER_REC_T_CONF_DIN_2	(`BASE_OFFSET+'h0C08)
`define FRER_REC_T_CONF_DIN_3	(`BASE_OFFSET+'h0C0A)
`define FRER_REC_T_CONF_DIN_4	(`BASE_OFFSET+'h0C0C)
`define FRER_REC_T_CONF_DIN_5	(`BASE_OFFSET+'h0C0E)
`define FRER_REC_T_CONF_DIN_6	(`BASE_OFFSET+'h0C10)
`define FRER_REC_T_CONF_DIN_7	(`BASE_OFFSET+'h0C12)
`define FRER_REC_T_CONF_DIN_8	(`BASE_OFFSET+'h0C14)
`define FRER_REC_T_CONF_DOUT_0	(`BASE_OFFSET+'h0C16)
`define FRER_REC_T_CONF_DOUT_1	(`BASE_OFFSET+'h0C18)
`define FRER_REC_T_CONF_DOUT_2	(`BASE_OFFSET+'h0C1A)
`define FRER_REC_T_CONF_DOUT_3	(`BASE_OFFSET+'h0C1C)
`define FRER_REC_T_CONF_DOUT_4	(`BASE_OFFSET+'h0C1E)
`define FRER_REC_T_CONF_DOUT_5	(`BASE_OFFSET+'h0C20)
`define FRER_REC_T_CONF_DOUT_6	(`BASE_OFFSET+'h0C22)
`define FRER_REC_T_CONF_DOUT_7	(`BASE_OFFSET+'h0C24)
`define FRER_REC_T_CONF_DOUT_8	(`BASE_OFFSET+'h0C26)
`define FRER_AGE_TIMER	        (`BASE_OFFSET+'h0C2A)
`define RTAG_ETYPE	            (`BASE_OFFSET+'h0C40)
`define FRER_REC_DROP_R_TRIG	(`BASE_OFFSET+'h0C42)	
`define FRER_REC_DROP_ROUT_H	(`BASE_OFFSET+'h0C44)	
`define FRER_REC_DROP_ROUT_L	(`BASE_OFFSET+'h0C46)	
//`define RX_PTP_FORWARD_TABLE	
`define RX_PTP_FORWARD_TABLE_STATUS	    (`BASE_OFFSET+'h0E00)
`define RX_PTP_FORWARD_TABLE_CONTROL	(`BASE_OFFSET+'h0E02)	
`define RX_PTP_FORWARD_T_CONF_DIN_0	    (`BASE_OFFSET+'h0E04)	
`define RX_PTP_FORWARD_T_CONF_DIN_1	    (`BASE_OFFSET+'h0E06)
`define RX_PTP_FORWARD_T_CONF_DIN_2	    (`BASE_OFFSET+'h0E08)
`define RX_PTP_FORWARD_T_CONF_DOUT_0	(`BASE_OFFSET+'h0E0A)	
`define RX_PTP_FORWARD_T_CONF_DOUT_1	(`BASE_OFFSET+'h0E0C)
`define RX_PTP_FORWARD_T_CONF_DOUT_2	(`BASE_OFFSET+'h0E0E)	
`define CPU_PORT_CFG	(`BASE_OFFSET+'h0E20)	
`define HWE_PORT_CFG	(`BASE_OFFSET+'h0E22)	
// OUT_FP_TABLE	
`define OUT_FP_TABLE_STATUS	    (`BASE_OFFSET+'h1000)
`define OUT_FP_TABLE_CONTROL	(`BASE_OFFSET+'h1002)	
`define OUT_FP_T_CONF_DIN_0	    (`BASE_OFFSET+'h1004)	
`define OUT_FP_T_CONF_DIN_1	    (`BASE_OFFSET+'h1006)
`define OUT_FP_T_CONF_DIN_2	    (`BASE_OFFSET+'h1008)
`define OUT_FP_T_CONF_DIN_3	    (`BASE_OFFSET+'h100A)
`define OUT_FP_T_CONF_DIN_4	    (`BASE_OFFSET+'h100C)
`define OUT_FP_T_CONF_DOUT_0	(`BASE_OFFSET+'h100E)	
`define OUT_FP_T_CONF_DOUT_1	(`BASE_OFFSET+'h1010)
`define OUT_FP_T_CONF_DOUT_2	(`BASE_OFFSET+'h1012)
`define OUT_FP_T_CONF_DOUT_3	(`BASE_OFFSET+'h1014)
`define OUT_FP_T_CONF_DOUT_4	(`BASE_OFFSET+'h1016)
// L2_MC_TABLE	
`define L2_MC_TABLE_STATUS	(`BASE_OFFSET+'h1020)
`define L2_MC_TABLE_CONTROL	(`BASE_OFFSET+'h1022)
`define L2_MC_T_CONF_DIN_0	(`BASE_OFFSET+'h1024)	
`define L2_MC_T_CONF_DIN_1	(`BASE_OFFSET+'h1026)
`define L2_MC_T_CONF_DIN_2	(`BASE_OFFSET+'h1028)
`define L2_MC_T_CONF_DOUT_0	(`BASE_OFFSET+'h102A)	
`define L2_MC_T_CONF_DOUT_1	(`BASE_OFFSET+'h102C)
`define L2_MC_T_CONF_DOUT_2	(`BASE_OFFSET+'h102E)
`define RX_BC_DROP_R_TRIG	(`BASE_OFFSET+'h1040)
`define RX_BC_DROP_ROUT_H	(`BASE_OFFSET+'h1042)
`define RX_BC_DROP_ROUT_L	(`BASE_OFFSET+'h1044)
`define RX_UC_DROP_R_TRIG	(`BASE_OFFSET+'h1046)	
`define RX_UC_DROP_ROUT_H	(`BASE_OFFSET+'h1048)	
`define RX_UC_DROP_ROUT_L	(`BASE_OFFSET+'h104A)
`define RX_KMC_DROP_R_TRIG	(`BASE_OFFSET+'h104C)	
`define RX_KMC_DROP_ROUT_H	(`BASE_OFFSET+'h104E)
`define RX_KMC_DROP_ROUT_L	(`BASE_OFFSET+'h1050)
`define RX_UMC_DROP_R_TRIG	(`BASE_OFFSET+'h1052)	
`define RX_UMC_DROP_ROUT_H	(`BASE_OFFSET+'h1054)	
`define RX_UMC_DROP_ROUT_L	(`BASE_OFFSET+'h1056)
`define RX_DVP_DROP_R_TRIG	(`BASE_OFFSET+'h1058)	
`define RX_DVP_DROP_ROUT_H	(`BASE_OFFSET+'h105A)	
`define RX_DVP_DROP_ROUT_L	(`BASE_OFFSET+'h105C)

//EVLAN_XLATE_TABLE	
`define EVLAN_XLATE_TABLE_STATUS	(`BASE_OFFSET+'h0020)
`define EVLAN_XLATE_TABLE_CONTROL	(`BASE_OFFSET+'h0022)
`define EVLAN_XLATE_T_CONF_KEY	    (`BASE_OFFSET+'h0024)
`define EVLAN_XLATE_T_DIN_0	        (`BASE_OFFSET+'h0026)
`define EVLAN_XLATE_T_DIN_1	        (`BASE_OFFSET+'h0028)
`define EVLAN_XLATE_T_DOUT_0	    (`BASE_OFFSET+'h002A)
`define EVLAN_XLATE_T_DOUT_1	    (`BASE_OFFSET+'h002C)
`define EVLAN_XLATE_T_DOUT_2	    (`BASE_OFFSET+'h002E)	
// EVLAN_ACTION_TABLE	
`define EVLAN_ACTION_TABLE_STATUS	(`BASE_OFFSET+'h0040)
`define EVLAN_ACTION_TABLE_CONTROL	(`BASE_OFFSET+'h0042)
`define EVLAN_ACTION_T_CONF_DIN_0	(`BASE_OFFSET+'h0044)	
`define EVLAN_ACTION_T_CONF_DIN_1	(`BASE_OFFSET+'h0046)
`define EVLAN_ACTION_T_CONF_DOUT_0	(`BASE_OFFSET+'h0048)	
`define EVLAN_ACTION_T_CONF_DOUT_1	(`BASE_OFFSET+'h004A)
//`define EVLAN_PROPERTY_TABLE	
`define EVLAN_PROPERTY_TABLE_STATUS  	(`BASE_OFFSET+'h0060)
`define EVLAN_PROPERTY_TABLE_CONTROL	(`BASE_OFFSET+'h0062)
`define EVLAN_PROPERTY_T_CONF_DIN_0	    (`BASE_OFFSET+'h0064)	
`define EVLAN_PROPERTY_T_CONF_DIN_1	    (`BASE_OFFSET+'h0066)
`define EVLAN_PROPERTY_T_CONF_DIN_2	    (`BASE_OFFSET+'h0068)
`define EVLAN_PROPERTY_T_CONF_DIN_3	    (`BASE_OFFSET+'h006A)
`define EVLAN_PROPERTY_T_CONF_DOUT_0	(`BASE_OFFSET+'h006C)	
`define EVLAN_PROPERTY_T_CONF_DOUT_1	(`BASE_OFFSET+'h006E)
`define EVLAN_PROPERTY_T_CONF_DOUT_2	(`BASE_OFFSET+'h0070)
`define EVLAN_PROPERTY_T_CONF_DOUT_3	(`BASE_OFFSET+'h0072)	
// EVLAN_STG_TABLE	
`define EVLAN_STG_TABLE_STATUS	(`BASE_OFFSET+'h0080)
`define EVLAN_STG_TABLE_CONTROL	(`BASE_OFFSET+'h0082)
`define ESTG_T_CONF_DIN_0	    (`BASE_OFFSET+'h0084)
`define ESTG_T_CONF_DIN_1	    (`BASE_OFFSET+'h0086)
`define ESTG_T_CONF_DIN_2	    (`BASE_OFFSET+'h0088)
`define ESTG_T_CONF_DIN_3	    (`BASE_OFFSET+'h008A)
`define ESTG_T_CONF_DOUT_0	    (`BASE_OFFSET+'h008C)
`define ESTG_T_CONF_DOUT_1	    (`BASE_OFFSET+'h008E)
`define ESTG_T_CONF_DOUT_2	    (`BASE_OFFSET+'h0090)
`define ESTG_T_CONF_DOUT_3	    (`BASE_OFFSET+'h0092)	
`define EPP_IN_DROP_R_TRIG	    (`BASE_OFFSET+'h00A0)	
`define EPP_IN_DROP_ROUT_H	    (`BASE_OFFSET+'h00A2)	
`define EPP_IN_DROP_ROUT_L	    (`BASE_OFFSET+'h00A4)
`define STP_OUT_DROP_R_TRIG	    (`BASE_OFFSET+'h00A6)	
`define STP_OUT_DROP_ROUT_H	    (`BASE_OFFSET+'h00A8)	
`define STP_OUT_DROP_ROUT_L	    (`BASE_OFFSET+'h00AA)
// OPORT_PRO_TABLE	
`define OPORT_PRO_TABLE_STATUS	(`BASE_OFFSET+'h0200)
`define OPORT_PRO_TABLE_CONTROL	(`BASE_OFFSET+'h0202)
`define OPORT_PRO_TABLE_DIN_0	(`BASE_OFFSET+'h0204)	
`define OPORT_PRO_TABLE_DIN_1	(`BASE_OFFSET+'h0206)
`define OPORT_PRO_TABLE_DOUT_0	(`BASE_OFFSET+'h0208)	
`define OPORT_PRO_TABLE_DOUT_1	(`BASE_OFFSET+'h020A)
// DOT1P_MAP_TABLE	
`define DOT1P_MAP_TABLE_STATUS	(`BASE_OFFSET+'h0220)
`define DOT1P_MAP_TABLE_CONTROL	(`BASE_OFFSET+'h0222)
`define DOT1P_MAP_T_DIN_0	    (`BASE_OFFSET+'h0224)	
`define DOT1P_MAP_T_DIN_1	    (`BASE_OFFSET+'h0226)
`define DOT1P_MAP_T_DOUT_0	    (`BASE_OFFSET+'h0228)	
`define DOT1P_MAP_T_DOUT_1	    (`BASE_OFFSET+'h022a)	
// LAG_SEL_PORT_TABLE	
`define LAG_SEL_PORT_TABLE_STATUS	(`BASE_OFFSET+'h0240)
`define LAG_SEL_PORT_TABLE_CONTROL	(`BASE_OFFSET+'h0242)
`define LAG_SEL_PORT_T_CONF_DIN_0	(`BASE_OFFSET+'h0244)	
`define LAG_SEL_PORT_T_CONF_DIN_1	(`BASE_OFFSET+'h0246)
`define LAG_SEL_PORT_T_CONF_DOUT_0	(`BASE_OFFSET+'h0248)	
`define LAG_SEL_PORT_T_CONF_DOUT_1	(`BASE_OFFSET+'h024A)	
// O_PHY_PORT_PRO_TABLE	
`define O_PHY_PORT_PRO_TABLE_STATUS	    (`BASE_OFFSET+'h0260)
`define O_PHY_PORT_PRO_TABLE_CONTROL	(`BASE_OFFSET+'h0262)
`define O_PHY_PORT_PRO_T_CONF_DIN_0	    (`BASE_OFFSET+'h0264)	
`define O_PHY_PORT_PRO_T_CONF_DIN_1	    (`BASE_OFFSET+'h0266)
`define O_PHY_PORT_PRO_T_CONF_DIN_2	    (`BASE_OFFSET+'h0268)
`define O_PHY_PORT_PRO_T_CONF_DIN_3	    (`BASE_OFFSET+'h026A)
`define O_PHY_PORT_PRO_T_CONF_DIN_4	    (`BASE_OFFSET+'h026C)
`define O_PHY_PORT_PRO_T_CONF_DIN_5	    (`BASE_OFFSET+'h026E)
`define O_PHY_PORT_PRO_T_CONF_DIN_6	    (`BASE_OFFSET+'h0270)
`define O_PHY_PORT_PRO_T_CONF_DIN_7	    (`BASE_OFFSET+'h0272)
`define O_PHY_PORT_PRO_T_CONF_DOUT_0	(`BASE_OFFSET+'h0274)	
`define O_PHY_PORT_PRO_T_CONF_DOUT_1	(`BASE_OFFSET+'h0276)
`define O_PHY_PORT_PRO_T_CONF_DOUT_2	(`BASE_OFFSET+'h0278)
`define O_PHY_PORT_PRO_T_CONF_DOUT_3	(`BASE_OFFSET+'h027A)
`define O_PHY_PORT_PRO_T_CONF_DOUT_4	(`BASE_OFFSET+'h027C)
`define O_PHY_PORT_PRO_T_CONF_DOUT_5	(`BASE_OFFSET+'h027E)
`define O_PHY_PORT_PRO_T_CONF_DOUT_6	(`BASE_OFFSET+'h0280)
`define O_PHY_PORT_PRO_T_CONF_DOUT_7	(`BASE_OFFSET+'h0282)	
`define E_FILTER_DROP_R_TRIG	        (`BASE_OFFSET+'h02A0)	
`define IP_BIND_DROP_ROUT_H	            (`BASE_OFFSET+'h02A2)	
`define IP_BIND_DROP_ROUT_L	            (`BASE_OFFSET+'h02A4)

`define PORT_POLLING_WEIGHT_TABLE_CFG_TRIGGER	(`BASE_OFFSET_GATHER+'h000)
`define PORT_POLLING_WEIGHT_TABLE_CFG_ADDR	    (`BASE_OFFSET_GATHER+'h001)
`define PORT_POLLING_WEIGHT_TABLE_CFG_PORT_ID	(`BASE_OFFSET_GATHER+'h002)
`define PORT_POLLING_WEIGHT_TABLE_LOOKUP_DATA	(`BASE_OFFSET_GATHER+'h003)

