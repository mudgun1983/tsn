package obm_mac_dec;
	parameter OBM_MAC_BP = 4;
endpackage:obm_mac_dec
