//FILE_HEADER-------------------------------------------------------
// ZTE  Copyright  (c)
// ZTE Company Confidential
//------------------------------------------------------------------
// Project Name : ZXLTE xxxx
// FILE NAME    : serdes_channel_ipcore.v
// AUTHOR       : pi qiang
// Department   : ZTE-BBU System Dept
// Email        : pi.qiang@zte.com.cn
//------------------------------------------------------------------
// Module Hiberarchy:
//x             |----xxx1
//x             |----xxx2
//x xxx_xxx-----|----xxx3 (Ϊ��ģ���������һ����ģ��������û���²�ģ�飬�ɲ���)
//x             |----xxx4
//x             |----xxx5
//-----------------------------------------------------------------
// Release History:
//-----------------------------------------------------------------
// Version      Date      Author    Description
// 1.0        2016-4-25   piqiang   ԭʼ�汾˵����
//-----------------------------------------------------------------
// Main Function:(Describing main function of the module)
// a)xxxxxxxx
// b)xxxxxxxx
//-----------------------------------------------------------------
//REUSE ISSUES: xxxxxxxx          
//Reset Strategy: xxxxxxxx
//Clock Strategy: xxxxxxxx
//Critical Timing: xxxxxxxx
//Asynchronous Interface: xxxxxxxx
//END_HEADER-------------------------------------------------------- 

`timescale 1ps/1ps
module serdes_channel_ipcore #
  (
  parameter C_GT_TYPE                           =     "GTYE3" 
  )                    
  ( 
  //CPLL                    
  input  wire    [0:0]                          CHANNEL_GTNORTHREFCLK0            ,
  input  wire    [0:0]                          CHANNEL_GTNORTHREFCLK1            ,
  input  wire    [0:0]                          CHANNEL_GTREFCLK0                 ,
  input  wire    [0:0]                          CHANNEL_GTREFCLK1                 ,
  input  wire    [0:0]                          CHANNEL_GTSOUTHREFCLK0            ,
  input  wire    [0:0]                          CHANNEL_GTSOUTHREFCLK1            ,
  input  wire    [0:0]                          CHANNEL_CPLLRESET                 ,
  input  wire    [0:0]                          CHANNEL_CPLLPD                    ,
  input  wire    [0:0]                          CHANNEL_CPLLLOCKDETCLK            ,
  input  wire    [2:0]                          CHANNEL_CPLLREFCLKSEL             ,
  output wire    [0:0]                          CHANNEL_CPLLFBCLKLOST             ,
  output wire    [0:0]                          CHANNEL_CPLLREFCLKLOST            ,
  output wire    [0:0]                          CHANNEL_CPLLLOCK                  ,
  //FROM QPLL
  input  wire    [0:0]                          CHANNEL_QPLL0CLK                  ,
  input  wire    [0:0]                          CHANNEL_QPLL0REFCLK               ,
  input  wire    [0:0]                          CHANNEL_QPLL1CLK                  ,
  input  wire    [0:0]                          CHANNEL_QPLL1REFCLK               ,
  //DRP
  input  wire    [0:0]                          CHANNEL_DRPCLK                    ,
  input  wire    [9:0]                          CHANNEL_DRPADDR                   ,
  input  wire    [15:0]                         CHANNEL_DRPDI                     ,
  input  wire    [0:0]                          CHANNEL_DRPWE                     ,
  input  wire    [0:0]                          CHANNEL_DRPEN                     ,
  output wire    [15:0]                         CHANNEL_DRPDO                     ,
  output wire    [0:0]                          CHANNEL_DRPRDY                    ,
  //   
  input  wire    [2:0]                          CHANNEL_LOOPBACK                  ,
  output wire    [0:0]                          CHANNEL_GTPOWERGOOD               ,
  //TX CLK
  input  wire    [1:0]                          CHANNEL_TXPLLCLKSEL               ,
  input  wire    [1:0]                          CHANNEL_TXSYSCLKSEL               ,
  input  wire    [2:0]                          CHANNEL_TXOUTCLKSEL               ,
  input  wire    [0:0]                          CHANNEL_TXPROGDIVRESET            ,
  output wire    [0:0]                          CHANNEL_TXPRGDIVRESETDONE         ,
  output wire    [0:0]                          CHANNEL_TXOUTCLK                  ,
  input  wire    [0:0]                          CHANNEL_TXUSRCLK                  ,
  input  wire    [0:0]                          CHANNEL_TXUSRCLK2                 ,
  //TX INTERFACE DATA
  input  wire    [7:0]                          CHANNEL_TXCTRL2                   ,
  input  wire    [127:0]                        CHANNEL_TXDATA                    ,
  //TX GEARBOX
  input  wire    [6:0]                          CHANNEL_TXSEQUENCE                ,
  input  wire    [5:0]                          CHANNEL_TXHEADER                  ,
  //TX 8B10B
  input  wire    [0:0]                          CHANNEL_TX8B10BEN                 ,
  //TX PRBS
  input  wire    [0:0]                          CHANNEL_TXPRBSFORCEERR            ,
  input  wire    [3:0]                          CHANNEL_TXPRBSSEL                 ,
  //TX BUFFER     
  output wire    [1:0]                          CHANNEL_TXBUFSTATUS               ,
  //TX Configurable Driver
  input  wire    [4:0]                          CHANNEL_TXDIFFCTRL                ,
  input  wire    [4:0]                          CHANNEL_TXPOSTCURSOR              ,
  input  wire    [4:0]                          CHANNEL_TXPRECURSOR               ,
  input  wire    [0:0]                          CHANNEL_TXINHIBIT                 ,
  //TX PIN DATA
  output wire    [0:0]                          CHANNEL_GTTXN                     ,
  output wire    [0:0]                          CHANNEL_GTTXP                     ,
  //TX OTHER                  
  input  wire    [1:0]                          CHANNEL_TXPD                      ,
  input  wire    [0:0]                          CHANNEL_GTTXRESET                 ,
  input  wire    [0:0]                          CHANNEL_TXUSERRDY                 ,
  output wire    [0:0]                          CHANNEL_TXRESETDONE               ,
  output wire    [0:0]                          CHANNEL_TXPMARESETDONE            ,
  //RX CLK
  input  wire    [1:0]                          CHANNEL_RXPLLCLKSEL               ,
  input  wire    [1:0]                          CHANNEL_RXSYSCLKSEL               ,
  input  wire    [2:0]                          CHANNEL_RXOUTCLKSEL               ,
  input  wire    [0:0]                          CHANNEL_RXPROGDIVRESET            ,
  output wire    [0:0]                          CHANNEL_RXPRGDIVRESETDONE         ,
  output wire    [0:0]                          CHANNEL_RXOUTCLK                  ,
  input  wire    [0:0]                          CHANNEL_RXUSRCLK                  ,
  input  wire    [0:0]                          CHANNEL_RXUSRCLK2                 ,
  //RX PIN DATA
  input  wire    [0:0]                          CHANNEL_GTRXN                     ,
  input  wire    [0:0]                          CHANNEL_GTRXP                     ,
  //RX PMA
  input  wire    [0:0]                          CHANNEL_RXLPMEN                   ,
  input  wire    [0:0]                          CHANNEL_RXLPMHFHOLD               ,
  input  wire    [0:0]                          CHANNEL_RXLPMLFHOLD               ,
  input  wire    [0:0]                          CHANNEL_RXDFEAGCHOLD              ,
  input  wire    [0:0]                          CHANNEL_RXDFELFHOLD               ,
  output wire    [0:0]                          CHANNEL_RXCDRLOCK                 ,
  //RX PRBS
  input  wire    [0:0]                          CHANNEL_RXPRBSCNTRESET            ,
  input  wire    [3:0]                          CHANNEL_RXPRBSSEL                 ,
  output wire    [0:0]                          CHANNEL_RXPRBSERR                 ,
  //RX ALIGN                  
  input  wire    [0:0]                          CHANNEL_RXCOMMADETEN              ,
  input  wire    [0:0]                          CHANNEL_RXMCOMMAALIGNEN           ,
  input  wire    [0:0]                          CHANNEL_RXPCOMMAALIGNEN           ,
  output wire    [0:0]                          CHANNEL_RXBYTEISALIGNED           ,
  //RX 8B10B
  input  wire    [0:0]                          CHANNEL_RX8B10BEN                 ,
  output wire    [15:0]                         CHANNEL_RXCTRL1                   ,
  output wire    [7:0]                          CHANNEL_RXCTRL3                   ,
  //RX BUFFER
  output wire    [2:0]                          CHANNEL_RXBUFSTATUS               ,
  //RX GEARBOX
  input  wire    [0:0]                          CHANNEL_RXGEARBOXSLIP             ,
  output wire    [5:0]                          CHANNEL_RXHEADER                  ,
  output wire    [1:0]                          CHANNEL_RXHEADERVALID             ,
  //RX INTERFACE DATA
  output wire    [15:0]                         CHANNEL_RXCTRL0                   ,
  output wire    [127:0]                        CHANNEL_RXDATA                    ,
  //RX OTHER
  input  wire    [1:0]                          CHANNEL_RXPD                      ,
  input  wire    [0:0]                          CHANNEL_GTRXRESET                 ,
  input  wire    [0:0]                          CHANNEL_RXUSERRDY                 ,
  output wire    [0:0]                          CHANNEL_RXRESETDONE               ,
  output wire    [0:0]                          CHANNEL_RXPMARESETDONE           
);



generate 
    if (C_GT_TYPE == "GTYE4_25") //��ʼ����25G,��368.64M�ο�ʱ�ӵ�QPLL0
        begin : gen_serdes_gtye4_channel_wrapper_25
            serdes_gtye4_channel_wrapper_25     serdes_gtye4_channel_wrapper_25 
            (
            //inputs
            .GTYE4_CHANNEL_CDRSTEPDIR                     ( 1'H0                            ), 
            .GTYE4_CHANNEL_CDRSTEPSQ                      ( 1'H0                            ),
            .GTYE4_CHANNEL_CDRSTEPSX                      ( 1'H0                            ),
            .GTYE4_CHANNEL_CFGRESET                       ( 1'H0                            ),
            .GTYE4_CHANNEL_CLKRSVD0                       ( 1'H0                            ),
            .GTYE4_CHANNEL_CLKRSVD1                       ( 1'H0                            ),
            .GTYE4_CHANNEL_CPLLFREQLOCK                   ( 1'H0                            ),
            .GTYE4_CHANNEL_CPLLLOCKDETCLK                 ( CHANNEL_CPLLLOCKDETCLK          ),
            .GTYE4_CHANNEL_CPLLLOCKEN                     ( 1'H1                            ),
            .GTYE4_CHANNEL_CPLLPD                         ( CHANNEL_CPLLPD                  ),
            .GTYE4_CHANNEL_CPLLREFCLKSEL                  ( CHANNEL_CPLLREFCLKSEL           ),
            .GTYE4_CHANNEL_CPLLRESET                      ( CHANNEL_CPLLRESET               ),
            .GTYE4_CHANNEL_DMONFIFORESET                  ( 1'H0                            ),
            .GTYE4_CHANNEL_DMONITORCLK                    ( 1'H0                            ),
            .GTYE4_CHANNEL_DRPADDR                        ( CHANNEL_DRPADDR[9:0]            ),
            .GTYE4_CHANNEL_DRPCLK                         ( CHANNEL_DRPCLK                  ),
            .GTYE4_CHANNEL_DRPDI                          ( CHANNEL_DRPDI                   ),
            .GTYE4_CHANNEL_DRPEN                          ( CHANNEL_DRPEN                   ),
            .GTYE4_CHANNEL_DRPRST                         ( 1'H0                            ),
            .GTYE4_CHANNEL_DRPWE                          ( CHANNEL_DRPWE                   ),
            .GTYE4_CHANNEL_EYESCANRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_EYESCANTRIGGER                 ( 1'H0                            ),
            .GTYE4_CHANNEL_FREQOS                         ( 1'H0                            ),
            .GTYE4_CHANNEL_GTGREFCLK                      ( 1'H0                            ),
            .GTYE4_CHANNEL_GTNORTHREFCLK0                 ( CHANNEL_GTNORTHREFCLK0          ),
            .GTYE4_CHANNEL_GTNORTHREFCLK1                 ( CHANNEL_GTNORTHREFCLK1          ),
            .GTYE4_CHANNEL_GTREFCLK0                      ( CHANNEL_GTREFCLK0               ),
            .GTYE4_CHANNEL_GTREFCLK1                      ( CHANNEL_GTREFCLK1               ),
            .GTYE4_CHANNEL_GTRSVD                         ( 16'H0000                        ),
            .GTYE4_CHANNEL_GTRXRESET                      ( CHANNEL_GTRXRESET               ),
            .GTYE4_CHANNEL_GTRXRESETSEL                   ( 1'H0                            ),
            .GTYE4_CHANNEL_GTSOUTHREFCLK0                 ( CHANNEL_GTSOUTHREFCLK0          ),
            .GTYE4_CHANNEL_GTSOUTHREFCLK1                 ( CHANNEL_GTSOUTHREFCLK1          ),
            .GTYE4_CHANNEL_GTTXRESET                      ( CHANNEL_GTTXRESET               ),
            .GTYE4_CHANNEL_GTTXRESETSEL                   ( 1'H0                            ),
            .GTYE4_CHANNEL_GTYRXN                         ( CHANNEL_GTRXN                   ),
            .GTYE4_CHANNEL_GTYRXP                         ( CHANNEL_GTRXP                   ),
            .GTYE4_CHANNEL_INCPCTRL                       ( 1'H0                            ),
            .GTYE4_CHANNEL_LOOPBACK                       ( CHANNEL_LOOPBACK                ),
            .GTYE4_CHANNEL_PCIEEQRXEQADAPTDONE            ( 1'H0                            ),
            .GTYE4_CHANNEL_PCIERSTIDLE                    ( 1'H0                            ),
            .GTYE4_CHANNEL_PCIERSTTXSYNCSTART             ( 1'H0                            ),
            .GTYE4_CHANNEL_PCIEUSERRATEDONE               ( 1'H0                            ),
            .GTYE4_CHANNEL_PCSRSVDIN                      ( 16'H0000                        ),
            .GTYE4_CHANNEL_QPLL0CLK                       ( CHANNEL_QPLL0CLK                ),
            .GTYE4_CHANNEL_QPLL0FREQLOCK                  ( 1'H0                            ),
            .GTYE4_CHANNEL_QPLL0REFCLK                    ( CHANNEL_QPLL0REFCLK             ),
            .GTYE4_CHANNEL_QPLL1CLK                       ( CHANNEL_QPLL1CLK                ),
            .GTYE4_CHANNEL_QPLL1FREQLOCK                  ( 1'H0                            ),
            .GTYE4_CHANNEL_QPLL1REFCLK                    ( CHANNEL_QPLL1REFCLK             ),
            .GTYE4_CHANNEL_RESETOVRD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RX8B10BEN                      ( CHANNEL_RX8B10BEN               ),
            .GTYE4_CHANNEL_RXAFECFOKEN                    ( 1'H1                            ),
            .GTYE4_CHANNEL_RXBUFRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDRFREQRESET                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDRHOLD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDROVRDEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDRRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDEN                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDI                      ( 5'H00                           ),
            .GTYE4_CHANNEL_RXCHBONDLEVEL                  ( 3'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDMASTER                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDSLAVE                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCKCALRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCKCALSTART                   ( 7'H00                           ),
            .GTYE4_CHANNEL_RXCOMMADETEN                   ( CHANNEL_RXCOMMADETEN            ),
            .GTYE4_CHANNEL_RXDFEAGCHOLD                   ( CHANNEL_RXDFEAGCHOLD            ),
            .GTYE4_CHANNEL_RXDFEAGCOVRDEN                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKFCNUM                 ( 4'HD                            ),
            .GTYE4_CHANNEL_RXDFECFOKFEN                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKFPULSE                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKHOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKOVREN                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEKHHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEKHOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFELFHOLD                    ( CHANNEL_RXDFELFHOLD             ),
            .GTYE4_CHANNEL_RXDFELFOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFELPMRESET                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP10HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP10OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP11HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP11OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP12HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP12OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP13HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP13OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP14HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP14OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP15HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP15OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP2HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP2OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP3HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP3OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP4HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP4OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP5HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP5OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP6HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP6OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP7HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP7OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP8HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP8OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP9HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP9OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEUTHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEUTOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEVPHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEVPOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEXYDEN                     ( 1'H1                            ),
            .GTYE4_CHANNEL_RXDLYBYPASS                    ( 1'H1                            ),
            .GTYE4_CHANNEL_RXDLYEN                        ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDLYOVRDEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDLYSRESET                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXELECIDLEMODE                 ( 2'H3                            ),
            .GTYE4_CHANNEL_RXEQTRAINING                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXGEARBOXSLIP                  ( CHANNEL_RXGEARBOXSLIP           ),
            .GTYE4_CHANNEL_RXLATCLK                       ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMEN                        ( CHANNEL_RXLPMEN                 ),
            .GTYE4_CHANNEL_RXLPMGCHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMGCOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMHFHOLD                    ( CHANNEL_RXLPMHFHOLD             ),
            .GTYE4_CHANNEL_RXLPMHFOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMLFHOLD                    ( CHANNEL_RXLPMLFHOLD             ),
            .GTYE4_CHANNEL_RXLPMLFKLOVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMOSHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMOSOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXMCOMMAALIGNEN                ( CHANNEL_RXMCOMMAALIGNEN         ),
            .GTYE4_CHANNEL_RXMONITORSEL                   ( 2'H0                            ),
            .GTYE4_CHANNEL_RXOOBRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOSCALRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOSHOLD                       ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOSOVRDEN                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOUTCLKSEL                    ( CHANNEL_RXOUTCLKSEL             ),
            .GTYE4_CHANNEL_RXPCOMMAALIGNEN                ( CHANNEL_RXPCOMMAALIGNEN         ),
            .GTYE4_CHANNEL_RXPCSRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPD                           ( CHANNEL_RXPD                    ),
            .GTYE4_CHANNEL_RXPHALIGN                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPHALIGNEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPHDLYPD                      ( 1'H1                            ),
            .GTYE4_CHANNEL_RXPHDLYRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPLLCLKSEL                    ( CHANNEL_RXPLLCLKSEL             ),
            .GTYE4_CHANNEL_RXPMARESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPOLARITY                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPRBSCNTRESET                 ( CHANNEL_RXPRBSCNTRESET          ),
            .GTYE4_CHANNEL_RXPRBSSEL                      ( CHANNEL_RXPRBSSEL               ),
            .GTYE4_CHANNEL_RXPROGDIVRESET                 ( CHANNEL_RXPROGDIVRESET          ),
            .GTYE4_CHANNEL_RXRATE                         ( 3'H0                            ),
            .GTYE4_CHANNEL_RXRATEMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSLIDE                        ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSLIPOUTCLK                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSLIPPMA                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYNCALLIN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYNCIN                       ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYNCMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYSCLKSEL                    ( CHANNEL_RXSYSCLKSEL             ),
            .GTYE4_CHANNEL_RXTERMINATION                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXUSERRDY                      ( CHANNEL_RXUSERRDY               ),
            .GTYE4_CHANNEL_RXUSRCLK                       ( CHANNEL_RXUSRCLK                ),
            .GTYE4_CHANNEL_RXUSRCLK2                      ( CHANNEL_RXUSRCLK2               ),
            .GTYE4_CHANNEL_SIGVALIDCLK                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TSTIN                          ( 20'H00000                       ),
            .GTYE4_CHANNEL_TX8B10BBYPASS                  ( 8'H00                           ),
            .GTYE4_CHANNEL_TX8B10BEN                      ( CHANNEL_TX8B10BEN               ),
            .GTYE4_CHANNEL_TXCOMINIT                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXCOMSAS                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXCOMWAKE                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXCTRL0                        ( 16'H0000                        ),
            .GTYE4_CHANNEL_TXCTRL1                        ( 16'H0000                        ),
            .GTYE4_CHANNEL_TXCTRL2                        ( CHANNEL_TXCTRL2                 ),
            .GTYE4_CHANNEL_TXDATA                         ( CHANNEL_TXDATA                  ),
            .GTYE4_CHANNEL_TXDATAEXTENDRSVD               ( 8'H00                           ),
            .GTYE4_CHANNEL_TXDCCFORCESTART                ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDCCRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDEEMPH                       ( 2'H0                            ),
            .GTYE4_CHANNEL_TXDETECTRX                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDIFFCTRL                     ( CHANNEL_TXDIFFCTRL[4:0]         ),
            .GTYE4_CHANNEL_TXDLYBYPASS                    ( 1'H1                            ),
            .GTYE4_CHANNEL_TXDLYEN                        ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYHOLD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYOVRDEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYSRESET                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYUPDOWN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXELECIDLE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXHEADER                       ( CHANNEL_TXHEADER                ),
            .GTYE4_CHANNEL_TXINHIBIT                      ( CHANNEL_TXINHIBIT               ),
            .GTYE4_CHANNEL_TXLATCLK                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXLFPSTRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_TXLFPSU2LPEXIT                 ( 1'H0                            ),
            .GTYE4_CHANNEL_TXLFPSU3WAKE                   ( 1'H0                            ),
            .GTYE4_CHANNEL_TXMAINCURSOR                   ( 7'H00                           ),
            .GTYE4_CHANNEL_TXMARGIN                       ( 3'H0                            ),
            .GTYE4_CHANNEL_TXMUXDCDEXHOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_TXMUXDCDORWREN                 ( 1'H0                            ),
            .GTYE4_CHANNEL_TXONESZEROS                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXOUTCLKSEL                    ( CHANNEL_TXOUTCLKSEL             ),
            .GTYE4_CHANNEL_TXPCSRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPD                           ( CHANNEL_TXPD                    ),
            .GTYE4_CHANNEL_TXPDELECIDLEMODE               ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHALIGN                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHALIGNEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHDLYPD                      ( 1'H1                            ),
            .GTYE4_CHANNEL_TXPHDLYRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHDLYTSTCLK                  ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHINIT                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHOVRDEN                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMEN                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMPD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMSEL                     ( 1'H1                            ),
            .GTYE4_CHANNEL_TXPIPPMSTEPSIZE                ( 5'H00                           ),
            .GTYE4_CHANNEL_TXPISOPD                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPLLCLKSEL                    ( CHANNEL_TXPLLCLKSEL             ),
            .GTYE4_CHANNEL_TXPMARESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPOLARITY                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPOSTCURSOR                   ( CHANNEL_TXPOSTCURSOR            ),
            .GTYE4_CHANNEL_TXPRBSFORCEERR                 ( CHANNEL_TXPRBSFORCEERR          ),
            .GTYE4_CHANNEL_TXPRBSSEL                      ( CHANNEL_TXPRBSSEL               ),
            .GTYE4_CHANNEL_TXPRECURSOR                    ( CHANNEL_TXPRECURSOR             ),
            .GTYE4_CHANNEL_TXPROGDIVRESET                 ( CHANNEL_TXPROGDIVRESET          ),
            .GTYE4_CHANNEL_TXRATE                         ( 3'H0                            ),
            .GTYE4_CHANNEL_TXRATEMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSEQUENCE                     ( CHANNEL_TXSEQUENCE              ),
            .GTYE4_CHANNEL_TXSWING                        ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYNCALLIN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYNCIN                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYNCMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYSCLKSEL                    ( CHANNEL_TXSYSCLKSEL             ),
            .GTYE4_CHANNEL_TXUSERRDY                      ( CHANNEL_TXUSERRDY               ),
            .GTYE4_CHANNEL_TXUSRCLK                       ( CHANNEL_TXUSRCLK                ),
            .GTYE4_CHANNEL_TXUSRCLK2                      ( CHANNEL_TXUSRCLK2               ),
                                                           
            // outputs                                     
            .GTYE4_CHANNEL_BUFGTCE                        (                                 ),
            .GTYE4_CHANNEL_BUFGTCEMASK                    (                                 ),
            .GTYE4_CHANNEL_BUFGTDIV                       (                                 ),
            .GTYE4_CHANNEL_BUFGTRESET                     (                                 ),
            .GTYE4_CHANNEL_BUFGTRSTMASK                   (                                 ),
            .GTYE4_CHANNEL_CPLLFBCLKLOST                  ( CHANNEL_CPLLFBCLKLOST           ),
            .GTYE4_CHANNEL_CPLLLOCK                       ( CHANNEL_CPLLLOCK                ),
            .GTYE4_CHANNEL_CPLLREFCLKLOST                 ( CHANNEL_CPLLREFCLKLOST          ),
            .GTYE4_CHANNEL_DMONITOROUT                    (                                 ),
            .GTYE4_CHANNEL_DMONITOROUTCLK                 (                                 ),
            .GTYE4_CHANNEL_DRPDO                          ( CHANNEL_DRPDO                   ),
            .GTYE4_CHANNEL_DRPRDY                         ( CHANNEL_DRPRDY                  ),
            .GTYE4_CHANNEL_EYESCANDATAERROR               (                                 ),
            .GTYE4_CHANNEL_GTPOWERGOOD                    ( CHANNEL_GTPOWERGOOD             ),
            .GTYE4_CHANNEL_GTREFCLKMONITOR                (                                 ),
            .GTYE4_CHANNEL_GTYTXN                         ( CHANNEL_GTTXN                   ),
            .GTYE4_CHANNEL_GTYTXP                         ( CHANNEL_GTTXP                   ),
            .GTYE4_CHANNEL_PCIERATEGEN3                   (                                 ),
            .GTYE4_CHANNEL_PCIERATEIDLE                   (                                 ),
            .GTYE4_CHANNEL_PCIERATEQPLLPD                 (                                 ),
            .GTYE4_CHANNEL_PCIERATEQPLLRESET              (                                 ),
            .GTYE4_CHANNEL_PCIESYNCTXSYNCDONE             (                                 ),
            .GTYE4_CHANNEL_PCIEUSERGEN3RDY                (                                 ),
            .GTYE4_CHANNEL_PCIEUSERPHYSTATUSRST           (                                 ),
            .GTYE4_CHANNEL_PCIEUSERRATESTART              (                                 ),
            .GTYE4_CHANNEL_PCSRSVDOUT                     (                                 ),
            .GTYE4_CHANNEL_PHYSTATUS                      (                                 ),
            .GTYE4_CHANNEL_PINRSRVDAS                     (                                 ),
            .GTYE4_CHANNEL_POWERPRESENT                   (                                 ),
            .GTYE4_CHANNEL_RESETEXCEPTION                 (                                 ),
            .GTYE4_CHANNEL_RXBUFSTATUS                    ( CHANNEL_RXBUFSTATUS             ),
            .GTYE4_CHANNEL_RXBYTEISALIGNED                ( CHANNEL_RXBYTEISALIGNED         ),
            .GTYE4_CHANNEL_RXBYTEREALIGN                  (                                 ),
            .GTYE4_CHANNEL_RXCDRLOCK                      ( CHANNEL_RXCDRLOCK               ),
            .GTYE4_CHANNEL_RXCDRPHDONE                    (                                 ),
            .GTYE4_CHANNEL_RXCHANBONDSEQ                  (                                 ),
            .GTYE4_CHANNEL_RXCHANISALIGNED                (                                 ),
            .GTYE4_CHANNEL_RXCHANREALIGN                  (                                 ),
            .GTYE4_CHANNEL_RXCHBONDO                      (                                 ),
            .GTYE4_CHANNEL_RXCKCALDONE                    (                                 ),
            .GTYE4_CHANNEL_RXCLKCORCNT                    (                                 ),
            .GTYE4_CHANNEL_RXCOMINITDET                   (                                 ),
            .GTYE4_CHANNEL_RXCOMMADET                     (                                 ),
            .GTYE4_CHANNEL_RXCOMSASDET                    (                                 ),
            .GTYE4_CHANNEL_RXCOMWAKEDET                   (                                 ),
            .GTYE4_CHANNEL_RXCTRL0                        ( CHANNEL_RXCTRL0                 ),
            .GTYE4_CHANNEL_RXCTRL1                        ( CHANNEL_RXCTRL1                 ),
            .GTYE4_CHANNEL_RXCTRL2                        (                                 ),
            .GTYE4_CHANNEL_RXCTRL3                        ( CHANNEL_RXCTRL3                 ),
            .GTYE4_CHANNEL_RXDATA                         ( CHANNEL_RXDATA                  ),
            .GTYE4_CHANNEL_RXDATAEXTENDRSVD               (                                 ),
            .GTYE4_CHANNEL_RXDATAVALID                    (                                 ),
            .GTYE4_CHANNEL_RXDLYSRESETDONE                (                                 ),
            .GTYE4_CHANNEL_RXELECIDLE                     (                                 ),
            .GTYE4_CHANNEL_RXHEADER                       ( CHANNEL_RXHEADER                ),
            .GTYE4_CHANNEL_RXHEADERVALID                  ( CHANNEL_RXHEADERVALID           ),
            .GTYE4_CHANNEL_RXLFPSTRESETDET                (                                 ),
            .GTYE4_CHANNEL_RXLFPSU2LPEXITDET              (                                 ),
            .GTYE4_CHANNEL_RXLFPSU3WAKEDET                (                                 ),
            .GTYE4_CHANNEL_RXMONITOROUT                   (                                 ),
            .GTYE4_CHANNEL_RXOSINTDONE                    (                                 ),
            .GTYE4_CHANNEL_RXOSINTSTARTED                 (                                 ),
            .GTYE4_CHANNEL_RXOSINTSTROBEDONE              (                                 ),
            .GTYE4_CHANNEL_RXOSINTSTROBESTARTED           (                                 ),
            .GTYE4_CHANNEL_RXOUTCLK                       ( CHANNEL_RXOUTCLK                ),
            .GTYE4_CHANNEL_RXOUTCLKFABRIC                 (                                 ),
            .GTYE4_CHANNEL_RXOUTCLKPCS                    (                                 ),
            .GTYE4_CHANNEL_RXPHALIGNDONE                  (                                 ),
            .GTYE4_CHANNEL_RXPHALIGNERR                   (                                 ),
            .GTYE4_CHANNEL_RXPMARESETDONE                 ( CHANNEL_RXPMARESETDONE          ),
            .GTYE4_CHANNEL_RXPRBSERR                      ( CHANNEL_RXPRBSERR               ),
            .GTYE4_CHANNEL_RXPRBSLOCKED                   (                                 ),
            .GTYE4_CHANNEL_RXPRGDIVRESETDONE              ( CHANNEL_RXPRGDIVRESETDONE       ),
            .GTYE4_CHANNEL_RXRATEDONE                     (                                 ),
            .GTYE4_CHANNEL_RXRECCLKOUT                    (                                 ),
            .GTYE4_CHANNEL_RXRESETDONE                    ( CHANNEL_RXRESETDONE             ),
            .GTYE4_CHANNEL_RXSLIDERDY                     (                                 ),
            .GTYE4_CHANNEL_RXSLIPDONE                     (                                 ),
            .GTYE4_CHANNEL_RXSLIPOUTCLKRDY                (                                 ),
            .GTYE4_CHANNEL_RXSLIPPMARDY                   (                                 ),
            .GTYE4_CHANNEL_RXSTARTOFSEQ                   (                                 ),
            .GTYE4_CHANNEL_RXSTATUS                       (                                 ),
            .GTYE4_CHANNEL_RXSYNCDONE                     (                                 ),
            .GTYE4_CHANNEL_RXSYNCOUT                      (                                 ),
            .GTYE4_CHANNEL_RXVALID                        (                                 ),
            .GTYE4_CHANNEL_TXBUFSTATUS                    ( CHANNEL_TXBUFSTATUS             ),
            .GTYE4_CHANNEL_TXCOMFINISH                    (                                 ),
            .GTYE4_CHANNEL_TXDCCDONE                      (                                 ),
            .GTYE4_CHANNEL_TXDLYSRESETDONE                (                                 ),
            .GTYE4_CHANNEL_TXOUTCLK                       ( CHANNEL_TXOUTCLK                ),
            .GTYE4_CHANNEL_TXOUTCLKFABRIC                 (                                 ),
            .GTYE4_CHANNEL_TXOUTCLKPCS                    (                                 ),
            .GTYE4_CHANNEL_TXPHALIGNDONE                  (                                 ),
            .GTYE4_CHANNEL_TXPHINITDONE                   (                                 ),
            .GTYE4_CHANNEL_TXPMARESETDONE                 ( CHANNEL_TXPMARESETDONE          ),
            .GTYE4_CHANNEL_TXPRGDIVRESETDONE              ( CHANNEL_TXPRGDIVRESETDONE       ),
            .GTYE4_CHANNEL_TXRATEDONE                     (                                 ),
            .GTYE4_CHANNEL_TXRESETDONE                    ( CHANNEL_TXRESETDONE             ),
            .GTYE4_CHANNEL_TXSYNCDONE                     (                                 ),
            .GTYE4_CHANNEL_TXSYNCOUT                      (                                 )
            );
        end



    else if (C_GT_TYPE == "GTYE4_12") //��ʼ����12G,��368.64M�ο�ʱ�ӵ�QPLL0
        begin : gen_serdes_gtye4_channel_wrapper_12
            serdes_gtye4_channel_wrapper_12     serdes_gtye4_channel_wrapper_12 
            (
            //inputs
            .GTYE4_CHANNEL_CDRSTEPDIR                     ( 1'H0                            ), 
            .GTYE4_CHANNEL_CDRSTEPSQ                      ( 1'H0                            ),
            .GTYE4_CHANNEL_CDRSTEPSX                      ( 1'H0                            ),
            .GTYE4_CHANNEL_CFGRESET                       ( 1'H0                            ),
            .GTYE4_CHANNEL_CLKRSVD0                       ( 1'H0                            ),
            .GTYE4_CHANNEL_CLKRSVD1                       ( 1'H0                            ),
            .GTYE4_CHANNEL_CPLLFREQLOCK                   ( 1'H0                            ),
            .GTYE4_CHANNEL_CPLLLOCKDETCLK                 ( CHANNEL_CPLLLOCKDETCLK          ),
            .GTYE4_CHANNEL_CPLLLOCKEN                     ( 1'H1                            ),
            .GTYE4_CHANNEL_CPLLPD                         ( CHANNEL_CPLLPD                  ),
            .GTYE4_CHANNEL_CPLLREFCLKSEL                  ( CHANNEL_CPLLREFCLKSEL           ),
            .GTYE4_CHANNEL_CPLLRESET                      ( CHANNEL_CPLLRESET               ),
            .GTYE4_CHANNEL_DMONFIFORESET                  ( 1'H0                            ),
            .GTYE4_CHANNEL_DMONITORCLK                    ( 1'H0                            ),
            .GTYE4_CHANNEL_DRPADDR                        ( CHANNEL_DRPADDR[9:0]            ),
            .GTYE4_CHANNEL_DRPCLK                         ( CHANNEL_DRPCLK                  ),
            .GTYE4_CHANNEL_DRPDI                          ( CHANNEL_DRPDI                   ),
            .GTYE4_CHANNEL_DRPEN                          ( CHANNEL_DRPEN                   ),
            .GTYE4_CHANNEL_DRPRST                         ( 1'H0                            ),
            .GTYE4_CHANNEL_DRPWE                          ( CHANNEL_DRPWE                   ),
            .GTYE4_CHANNEL_EYESCANRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_EYESCANTRIGGER                 ( 1'H0                            ),
            .GTYE4_CHANNEL_FREQOS                         ( 1'H0                            ),
            .GTYE4_CHANNEL_GTGREFCLK                      ( 1'H0                            ),
            .GTYE4_CHANNEL_GTNORTHREFCLK0                 ( CHANNEL_GTNORTHREFCLK0          ),
            .GTYE4_CHANNEL_GTNORTHREFCLK1                 ( CHANNEL_GTNORTHREFCLK1          ),
            .GTYE4_CHANNEL_GTREFCLK0                      ( CHANNEL_GTREFCLK0               ),
            .GTYE4_CHANNEL_GTREFCLK1                      ( CHANNEL_GTREFCLK1               ),
            .GTYE4_CHANNEL_GTRSVD                         ( 16'H0000                        ),
            .GTYE4_CHANNEL_GTRXRESET                      ( CHANNEL_GTRXRESET               ),
            .GTYE4_CHANNEL_GTRXRESETSEL                   ( 1'H0                            ),
            .GTYE4_CHANNEL_GTSOUTHREFCLK0                 ( CHANNEL_GTSOUTHREFCLK0          ),
            .GTYE4_CHANNEL_GTSOUTHREFCLK1                 ( CHANNEL_GTSOUTHREFCLK1          ),
            .GTYE4_CHANNEL_GTTXRESET                      ( CHANNEL_GTTXRESET               ),
            .GTYE4_CHANNEL_GTTXRESETSEL                   ( 1'H0                            ),
            .GTYE4_CHANNEL_GTYRXN                         ( CHANNEL_GTRXN                   ),
            .GTYE4_CHANNEL_GTYRXP                         ( CHANNEL_GTRXP                   ),
            .GTYE4_CHANNEL_INCPCTRL                       ( 1'H0                            ),
            .GTYE4_CHANNEL_LOOPBACK                       ( CHANNEL_LOOPBACK                ),
            .GTYE4_CHANNEL_PCIEEQRXEQADAPTDONE            ( 1'H0                            ),
            .GTYE4_CHANNEL_PCIERSTIDLE                    ( 1'H0                            ),
            .GTYE4_CHANNEL_PCIERSTTXSYNCSTART             ( 1'H0                            ),
            .GTYE4_CHANNEL_PCIEUSERRATEDONE               ( 1'H0                            ),
            .GTYE4_CHANNEL_PCSRSVDIN                      ( 16'H0000                        ),
            .GTYE4_CHANNEL_QPLL0CLK                       ( CHANNEL_QPLL0CLK                ),
            .GTYE4_CHANNEL_QPLL0FREQLOCK                  ( 1'H0                            ),
            .GTYE4_CHANNEL_QPLL0REFCLK                    ( CHANNEL_QPLL0REFCLK             ),
            .GTYE4_CHANNEL_QPLL1CLK                       ( CHANNEL_QPLL1CLK                ),
            .GTYE4_CHANNEL_QPLL1FREQLOCK                  ( 1'H0                            ),
            .GTYE4_CHANNEL_QPLL1REFCLK                    ( CHANNEL_QPLL1REFCLK             ),
            .GTYE4_CHANNEL_RESETOVRD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RX8B10BEN                      ( CHANNEL_RX8B10BEN               ),
            .GTYE4_CHANNEL_RXAFECFOKEN                    ( 1'H1                            ),
            .GTYE4_CHANNEL_RXBUFRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDRFREQRESET                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDRHOLD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDROVRDEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCDRRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDEN                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDI                      ( 5'H00                           ),
            .GTYE4_CHANNEL_RXCHBONDLEVEL                  ( 3'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDMASTER                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCHBONDSLAVE                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCKCALRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXCKCALSTART                   ( 7'H00                           ),
            .GTYE4_CHANNEL_RXCOMMADETEN                   ( CHANNEL_RXCOMMADETEN            ),
            .GTYE4_CHANNEL_RXDFEAGCHOLD                   ( CHANNEL_RXDFEAGCHOLD            ),
            .GTYE4_CHANNEL_RXDFEAGCOVRDEN                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKFCNUM                 ( 4'HD                            ),
            .GTYE4_CHANNEL_RXDFECFOKFEN                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKFPULSE                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKHOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFECFOKOVREN                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEKHHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEKHOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFELFHOLD                    ( CHANNEL_RXDFELFHOLD             ),
            .GTYE4_CHANNEL_RXDFELFOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFELPMRESET                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP10HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP10OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP11HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP11OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP12HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP12OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP13HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP13OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP14HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP14OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP15HOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP15OVRDEN               ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP2HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP2OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP3HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP3OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP4HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP4OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP5HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP5OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP6HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP6OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP7HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP7OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP8HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP8OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP9HOLD                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFETAP9OVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEUTHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEUTOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEVPHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEVPOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDFEXYDEN                     ( 1'H1                            ),
            .GTYE4_CHANNEL_RXDLYBYPASS                    ( 1'H1                            ),
            .GTYE4_CHANNEL_RXDLYEN                        ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDLYOVRDEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXDLYSRESET                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXELECIDLEMODE                 ( 2'H3                            ),
            .GTYE4_CHANNEL_RXEQTRAINING                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXGEARBOXSLIP                  ( CHANNEL_RXGEARBOXSLIP           ),
            .GTYE4_CHANNEL_RXLATCLK                       ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMEN                        ( CHANNEL_RXLPMEN                 ),
            .GTYE4_CHANNEL_RXLPMGCHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMGCOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMHFHOLD                    ( CHANNEL_RXLPMHFHOLD             ),
            .GTYE4_CHANNEL_RXLPMHFOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMLFHOLD                    ( CHANNEL_RXLPMLFHOLD             ),
            .GTYE4_CHANNEL_RXLPMLFKLOVRDEN                ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMOSHOLD                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXLPMOSOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXMCOMMAALIGNEN                ( CHANNEL_RXMCOMMAALIGNEN         ),
            .GTYE4_CHANNEL_RXMONITORSEL                   ( 2'H0                            ),
            .GTYE4_CHANNEL_RXOOBRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOSCALRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOSHOLD                       ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOSOVRDEN                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXOUTCLKSEL                    ( CHANNEL_RXOUTCLKSEL             ),
            .GTYE4_CHANNEL_RXPCOMMAALIGNEN                ( CHANNEL_RXPCOMMAALIGNEN         ),
            .GTYE4_CHANNEL_RXPCSRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPD                           ( CHANNEL_RXPD                    ),
            .GTYE4_CHANNEL_RXPHALIGN                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPHALIGNEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPHDLYPD                      ( 1'H1                            ),
            .GTYE4_CHANNEL_RXPHDLYRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPLLCLKSEL                    ( CHANNEL_RXPLLCLKSEL             ),
            .GTYE4_CHANNEL_RXPMARESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPOLARITY                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXPRBSCNTRESET                 ( CHANNEL_RXPRBSCNTRESET          ),
            .GTYE4_CHANNEL_RXPRBSSEL                      ( CHANNEL_RXPRBSSEL               ),
            .GTYE4_CHANNEL_RXPROGDIVRESET                 ( CHANNEL_RXPROGDIVRESET          ),
            .GTYE4_CHANNEL_RXRATE                         ( 3'H0                            ),
            .GTYE4_CHANNEL_RXRATEMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSLIDE                        ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSLIPOUTCLK                   ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSLIPPMA                      ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYNCALLIN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYNCIN                       ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYNCMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_RXSYSCLKSEL                    ( CHANNEL_RXSYSCLKSEL             ),
            .GTYE4_CHANNEL_RXTERMINATION                  ( 1'H0                            ),
            .GTYE4_CHANNEL_RXUSERRDY                      ( CHANNEL_RXUSERRDY               ),
            .GTYE4_CHANNEL_RXUSRCLK                       ( CHANNEL_RXUSRCLK                ),
            .GTYE4_CHANNEL_RXUSRCLK2                      ( CHANNEL_RXUSRCLK2               ),
            .GTYE4_CHANNEL_SIGVALIDCLK                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TSTIN                          ( 20'H00000                       ),
            .GTYE4_CHANNEL_TX8B10BBYPASS                  ( 8'H00                           ),
            .GTYE4_CHANNEL_TX8B10BEN                      ( CHANNEL_TX8B10BEN               ),
            .GTYE4_CHANNEL_TXCOMINIT                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXCOMSAS                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXCOMWAKE                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXCTRL0                        ( 16'H0000                        ),
            .GTYE4_CHANNEL_TXCTRL1                        ( 16'H0000                        ),
            .GTYE4_CHANNEL_TXCTRL2                        ( CHANNEL_TXCTRL2                 ),
            .GTYE4_CHANNEL_TXDATA                         ( CHANNEL_TXDATA                  ),
            .GTYE4_CHANNEL_TXDATAEXTENDRSVD               ( 8'H00                           ),
            .GTYE4_CHANNEL_TXDCCFORCESTART                ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDCCRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDEEMPH                       ( 2'H0                            ),
            .GTYE4_CHANNEL_TXDETECTRX                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDIFFCTRL                     ( CHANNEL_TXDIFFCTRL[4:0]         ),
            .GTYE4_CHANNEL_TXDLYBYPASS                    ( 1'H1                            ),
            .GTYE4_CHANNEL_TXDLYEN                        ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYHOLD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYOVRDEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYSRESET                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXDLYUPDOWN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXELECIDLE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXHEADER                       ( CHANNEL_TXHEADER                ),
            .GTYE4_CHANNEL_TXINHIBIT                      ( CHANNEL_TXINHIBIT               ),
            .GTYE4_CHANNEL_TXLATCLK                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXLFPSTRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_TXLFPSU2LPEXIT                 ( 1'H0                            ),
            .GTYE4_CHANNEL_TXLFPSU3WAKE                   ( 1'H0                            ),
            .GTYE4_CHANNEL_TXMAINCURSOR                   ( 7'H00                           ),
            .GTYE4_CHANNEL_TXMARGIN                       ( 3'H0                            ),
            .GTYE4_CHANNEL_TXMUXDCDEXHOLD                 ( 1'H0                            ),
            .GTYE4_CHANNEL_TXMUXDCDORWREN                 ( 1'H0                            ),
            .GTYE4_CHANNEL_TXONESZEROS                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXOUTCLKSEL                    ( CHANNEL_TXOUTCLKSEL             ),
            .GTYE4_CHANNEL_TXPCSRESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPD                           ( CHANNEL_TXPD                    ),
            .GTYE4_CHANNEL_TXPDELECIDLEMODE               ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHALIGN                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHALIGNEN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHDLYPD                      ( 1'H1                            ),
            .GTYE4_CHANNEL_TXPHDLYRESET                   ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHDLYTSTCLK                  ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHINIT                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPHOVRDEN                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMEN                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMOVRDEN                  ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMPD                      ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPIPPMSEL                     ( 1'H1                            ),
            .GTYE4_CHANNEL_TXPIPPMSTEPSIZE                ( 5'H00                           ),
            .GTYE4_CHANNEL_TXPISOPD                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPLLCLKSEL                    ( CHANNEL_TXPLLCLKSEL             ),
            .GTYE4_CHANNEL_TXPMARESET                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPOLARITY                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXPOSTCURSOR                   ( CHANNEL_TXPOSTCURSOR            ),
            .GTYE4_CHANNEL_TXPRBSFORCEERR                 ( CHANNEL_TXPRBSFORCEERR          ),
            .GTYE4_CHANNEL_TXPRBSSEL                      ( CHANNEL_TXPRBSSEL               ),
            .GTYE4_CHANNEL_TXPRECURSOR                    ( CHANNEL_TXPRECURSOR             ),
            .GTYE4_CHANNEL_TXPROGDIVRESET                 ( CHANNEL_TXPROGDIVRESET          ),
            .GTYE4_CHANNEL_TXRATE                         ( 3'H0                            ),
            .GTYE4_CHANNEL_TXRATEMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSEQUENCE                     ( CHANNEL_TXSEQUENCE              ),
            .GTYE4_CHANNEL_TXSWING                        ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYNCALLIN                    ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYNCIN                       ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYNCMODE                     ( 1'H0                            ),
            .GTYE4_CHANNEL_TXSYSCLKSEL                    ( CHANNEL_TXSYSCLKSEL             ),
            .GTYE4_CHANNEL_TXUSERRDY                      ( CHANNEL_TXUSERRDY               ),
            .GTYE4_CHANNEL_TXUSRCLK                       ( CHANNEL_TXUSRCLK                ),
            .GTYE4_CHANNEL_TXUSRCLK2                      ( CHANNEL_TXUSRCLK2               ),
                                                           
            // outputs                                     
            .GTYE4_CHANNEL_BUFGTCE                        (                                 ),
            .GTYE4_CHANNEL_BUFGTCEMASK                    (                                 ),
            .GTYE4_CHANNEL_BUFGTDIV                       (                                 ),
            .GTYE4_CHANNEL_BUFGTRESET                     (                                 ),
            .GTYE4_CHANNEL_BUFGTRSTMASK                   (                                 ),
            .GTYE4_CHANNEL_CPLLFBCLKLOST                  ( CHANNEL_CPLLFBCLKLOST           ),
            .GTYE4_CHANNEL_CPLLLOCK                       ( CHANNEL_CPLLLOCK                ),
            .GTYE4_CHANNEL_CPLLREFCLKLOST                 ( CHANNEL_CPLLREFCLKLOST          ),
            .GTYE4_CHANNEL_DMONITOROUT                    (                                 ),
            .GTYE4_CHANNEL_DMONITOROUTCLK                 (                                 ),
            .GTYE4_CHANNEL_DRPDO                          ( CHANNEL_DRPDO                   ),
            .GTYE4_CHANNEL_DRPRDY                         ( CHANNEL_DRPRDY                  ),
            .GTYE4_CHANNEL_EYESCANDATAERROR               (                                 ),
            .GTYE4_CHANNEL_GTPOWERGOOD                    ( CHANNEL_GTPOWERGOOD             ),
            .GTYE4_CHANNEL_GTREFCLKMONITOR                (                                 ),
            .GTYE4_CHANNEL_GTYTXN                         ( CHANNEL_GTTXN                   ),
            .GTYE4_CHANNEL_GTYTXP                         ( CHANNEL_GTTXP                   ),
            .GTYE4_CHANNEL_PCIERATEGEN3                   (                                 ),
            .GTYE4_CHANNEL_PCIERATEIDLE                   (                                 ),
            .GTYE4_CHANNEL_PCIERATEQPLLPD                 (                                 ),
            .GTYE4_CHANNEL_PCIERATEQPLLRESET              (                                 ),
            .GTYE4_CHANNEL_PCIESYNCTXSYNCDONE             (                                 ),
            .GTYE4_CHANNEL_PCIEUSERGEN3RDY                (                                 ),
            .GTYE4_CHANNEL_PCIEUSERPHYSTATUSRST           (                                 ),
            .GTYE4_CHANNEL_PCIEUSERRATESTART              (                                 ),
            .GTYE4_CHANNEL_PCSRSVDOUT                     (                                 ),
            .GTYE4_CHANNEL_PHYSTATUS                      (                                 ),
            .GTYE4_CHANNEL_PINRSRVDAS                     (                                 ),
            .GTYE4_CHANNEL_POWERPRESENT                   (                                 ),
            .GTYE4_CHANNEL_RESETEXCEPTION                 (                                 ),
            .GTYE4_CHANNEL_RXBUFSTATUS                    ( CHANNEL_RXBUFSTATUS             ),
            .GTYE4_CHANNEL_RXBYTEISALIGNED                ( CHANNEL_RXBYTEISALIGNED         ),
            .GTYE4_CHANNEL_RXBYTEREALIGN                  (                                 ),
            .GTYE4_CHANNEL_RXCDRLOCK                      ( CHANNEL_RXCDRLOCK               ),
            .GTYE4_CHANNEL_RXCDRPHDONE                    (                                 ),
            .GTYE4_CHANNEL_RXCHANBONDSEQ                  (                                 ),
            .GTYE4_CHANNEL_RXCHANISALIGNED                (                                 ),
            .GTYE4_CHANNEL_RXCHANREALIGN                  (                                 ),
            .GTYE4_CHANNEL_RXCHBONDO                      (                                 ),
            .GTYE4_CHANNEL_RXCKCALDONE                    (                                 ),
            .GTYE4_CHANNEL_RXCLKCORCNT                    (                                 ),
            .GTYE4_CHANNEL_RXCOMINITDET                   (                                 ),
            .GTYE4_CHANNEL_RXCOMMADET                     (                                 ),
            .GTYE4_CHANNEL_RXCOMSASDET                    (                                 ),
            .GTYE4_CHANNEL_RXCOMWAKEDET                   (                                 ),
            .GTYE4_CHANNEL_RXCTRL0                        ( CHANNEL_RXCTRL0                 ),
            .GTYE4_CHANNEL_RXCTRL1                        ( CHANNEL_RXCTRL1                 ),
            .GTYE4_CHANNEL_RXCTRL2                        (                                 ),
            .GTYE4_CHANNEL_RXCTRL3                        ( CHANNEL_RXCTRL3                 ),
            .GTYE4_CHANNEL_RXDATA                         ( CHANNEL_RXDATA                  ),
            .GTYE4_CHANNEL_RXDATAEXTENDRSVD               (                                 ),
            .GTYE4_CHANNEL_RXDATAVALID                    (                                 ),
            .GTYE4_CHANNEL_RXDLYSRESETDONE                (                                 ),
            .GTYE4_CHANNEL_RXELECIDLE                     (                                 ),
            .GTYE4_CHANNEL_RXHEADER                       ( CHANNEL_RXHEADER                ),
            .GTYE4_CHANNEL_RXHEADERVALID                  ( CHANNEL_RXHEADERVALID           ),
            .GTYE4_CHANNEL_RXLFPSTRESETDET                (                                 ),
            .GTYE4_CHANNEL_RXLFPSU2LPEXITDET              (                                 ),
            .GTYE4_CHANNEL_RXLFPSU3WAKEDET                (                                 ),
            .GTYE4_CHANNEL_RXMONITOROUT                   (                                 ),
            .GTYE4_CHANNEL_RXOSINTDONE                    (                                 ),
            .GTYE4_CHANNEL_RXOSINTSTARTED                 (                                 ),
            .GTYE4_CHANNEL_RXOSINTSTROBEDONE              (                                 ),
            .GTYE4_CHANNEL_RXOSINTSTROBESTARTED           (                                 ),
            .GTYE4_CHANNEL_RXOUTCLK                       ( CHANNEL_RXOUTCLK                ),
            .GTYE4_CHANNEL_RXOUTCLKFABRIC                 (                                 ),
            .GTYE4_CHANNEL_RXOUTCLKPCS                    (                                 ),
            .GTYE4_CHANNEL_RXPHALIGNDONE                  (                                 ),
            .GTYE4_CHANNEL_RXPHALIGNERR                   (                                 ),
            .GTYE4_CHANNEL_RXPMARESETDONE                 ( CHANNEL_RXPMARESETDONE          ),
            .GTYE4_CHANNEL_RXPRBSERR                      ( CHANNEL_RXPRBSERR               ),
            .GTYE4_CHANNEL_RXPRBSLOCKED                   (                                 ),
            .GTYE4_CHANNEL_RXPRGDIVRESETDONE              ( CHANNEL_RXPRGDIVRESETDONE       ),
            .GTYE4_CHANNEL_RXRATEDONE                     (                                 ),
            .GTYE4_CHANNEL_RXRECCLKOUT                    (                                 ),
            .GTYE4_CHANNEL_RXRESETDONE                    ( CHANNEL_RXRESETDONE             ),
            .GTYE4_CHANNEL_RXSLIDERDY                     (                                 ),
            .GTYE4_CHANNEL_RXSLIPDONE                     (                                 ),
            .GTYE4_CHANNEL_RXSLIPOUTCLKRDY                (                                 ),
            .GTYE4_CHANNEL_RXSLIPPMARDY                   (                                 ),
            .GTYE4_CHANNEL_RXSTARTOFSEQ                   (                                 ),
            .GTYE4_CHANNEL_RXSTATUS                       (                                 ),
            .GTYE4_CHANNEL_RXSYNCDONE                     (                                 ),
            .GTYE4_CHANNEL_RXSYNCOUT                      (                                 ),
            .GTYE4_CHANNEL_RXVALID                        (                                 ),
            .GTYE4_CHANNEL_TXBUFSTATUS                    ( CHANNEL_TXBUFSTATUS             ),
            .GTYE4_CHANNEL_TXCOMFINISH                    (                                 ),
            .GTYE4_CHANNEL_TXDCCDONE                      (                                 ),
            .GTYE4_CHANNEL_TXDLYSRESETDONE                (                                 ),
            .GTYE4_CHANNEL_TXOUTCLK                       ( CHANNEL_TXOUTCLK                ),
            .GTYE4_CHANNEL_TXOUTCLKFABRIC                 (                                 ),
            .GTYE4_CHANNEL_TXOUTCLKPCS                    (                                 ),
            .GTYE4_CHANNEL_TXPHALIGNDONE                  (                                 ),
            .GTYE4_CHANNEL_TXPHINITDONE                   (                                 ),
            .GTYE4_CHANNEL_TXPMARESETDONE                 ( CHANNEL_TXPMARESETDONE          ),
            .GTYE4_CHANNEL_TXPRGDIVRESETDONE              ( CHANNEL_TXPRGDIVRESETDONE       ),
            .GTYE4_CHANNEL_TXRATEDONE                     (                                 ),
            .GTYE4_CHANNEL_TXRESETDONE                    ( CHANNEL_TXRESETDONE             ),
            .GTYE4_CHANNEL_TXSYNCDONE                     (                                 ),
            .GTYE4_CHANNEL_TXSYNCOUT                      (                                 )
            );
        end






endgenerate        
        
endmodule

