library verilog;
use verilog.vl_types.all;
entity dcn_cpu_main is
    generic(
        VERSION_MONTH   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        VERSION_DAY     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        VERSION_HOUR    : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        VERSION_MINUTE  : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        reset           : in     vl_logic;
        sys_clk         : in     vl_logic;
        cpu_clk         : in     vl_logic;
        cpu_rst         : in     vl_logic;
        cpu_addr        : in     vl_logic_vector(7 downto 0);
        cpu_cs          : in     vl_logic;
        cpu_rd          : in     vl_logic;
        cpu_wr          : in     vl_logic;
        cpu_din         : in     vl_logic_vector(15 downto 0);
        cpu_dout        : out    vl_logic_vector(15 downto 0);
        vlan_to_shim0_tx: out    vl_logic_vector(15 downto 0);
        vlan_to_shim1_tx: out    vl_logic_vector(15 downto 0);
        vlan_to_shim0_rx: out    vl_logic_vector(15 downto 0);
        vlan_to_shim1_rx: out    vl_logic_vector(15 downto 0);
        packet_restore_fifo_rst_tx: out    vl_logic;
        packet_restore_fifo_rst_rx: out    vl_logic;
        shim_buf_fifo_rst: out    vl_logic;
        soft_tx_rst     : out    vl_logic;
        soft_rx_rst     : out    vl_logic;
        loop_en         : out    vl_logic_vector(2 downto 0);
        packet_gen_en   : out    vl_logic;
        tx_packet_rcv   : in     vl_logic;
        tx_crc_ind      : in     vl_logic;
        tx_packet_discard_shim0: in     vl_logic;
        tx_fifo_empty_shim0: in     vl_logic;
        tx_fifo_full_shim0: in     vl_logic;
        tx_fifo_data_cnt_shim0: in     vl_logic_vector(12 downto 0);
        tx_buf_fifo_empty_shim0: in     vl_logic;
        tx_buf_fifo_full_shim0: in     vl_logic;
        tx_packet_discard_shim1: in     vl_logic;
        tx_fifo_empty_shim1: in     vl_logic;
        tx_fifo_full_shim1: in     vl_logic;
        tx_fifo_data_cnt_shim1: in     vl_logic_vector(12 downto 0);
        tx_buf_fifo_empty_shim1: in     vl_logic;
        tx_buf_fifo_full_shim1: in     vl_logic;
        rx_packet_rcv   : in     vl_logic;
        rx_crc_ind      : in     vl_logic;
        rx_packet_discard_shim0: in     vl_logic;
        rx_fifo_empty_shim0: in     vl_logic;
        rx_fifo_full_shim0: in     vl_logic;
        rx_fifo_data_cnt_shim0: in     vl_logic_vector(12 downto 0);
        rx_packet_discard_shim1: in     vl_logic;
        rx_fifo_empty_shim1: in     vl_logic;
        rx_fifo_full_shim1: in     vl_logic;
        rx_fifo_data_cnt_shim1: in     vl_logic_vector(12 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of VERSION_MONTH : constant is 2;
    attribute mti_svvh_generic_type of VERSION_DAY : constant is 2;
    attribute mti_svvh_generic_type of VERSION_HOUR : constant is 2;
    attribute mti_svvh_generic_type of VERSION_MINUTE : constant is 2;
end dcn_cpu_main;
