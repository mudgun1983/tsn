library verilog;
use verilog.vl_types.all;
entity xgmii64_rx_if is
end xgmii64_rx_if;
