`include "src/obm_mac_interface.sv"
`include "src/obm_mac_dec.sv"
package obm_mac_package;
	import uvm_pkg::*;
	import base_package::*;
	`include "src/obm_mac_xaction.sv"
	`include "src/obm_mac_monitor.sv"
	`include "src/obm_mac_interface_agent.sv"
endpackage

import obm_mac_package::*;
