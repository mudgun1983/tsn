package crllist_chk_dec;
	parameter DATA_NS = 32'd1_000_000_000;
	parameter LAT_CYC_NUM  = 4;
	parameter CYC_PEROID   = 8;
	parameter GATE_LATENCY = (LAT_CYC_NUM*CYC_PEROID);
endpackage:crllist_chk_dec
