package base_package;
	import uvm_pkg::*;
	`include "./monitor_base.sv"
	`include "./component_base.sv"
	`include "./interface_agent_base.sv"
endpackage

import base_package::*;

