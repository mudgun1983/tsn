library verilog;
use verilog.vl_types.all;
entity cpu_pkg is
end cpu_pkg;
