`define U_SCATTER pcs_tb_top.UUT.tsn_sw_top.scatter
`define U_OBM(MAC_NUM) pcs_tb_top.UUT.tsn_sw_top.obm_top_``MAC_NUM``
