
class cpu_config extends uvm_object;

   `uvm_object_utils(cpu_config)
   virtual cpu_if vif;
  
endclass

