//PHY_PORT_TABLE
//`define DUMMY_DUT