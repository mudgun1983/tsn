library verilog;
use verilog.vl_types.all;
entity pcs_xilinx_serdes_if is
end pcs_xilinx_serdes_if;
