package obm_dut_cfg_package;
    import uvm_pkg::*;
	`include "obm_dut_cfg.sv"
	`include "obm_case0_cfg.sv"
endpackage

import obm_dut_cfg_package::*;
