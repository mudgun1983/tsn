`include "src/mac_tx_interface.sv"
package mac_tx_package;
	import uvm_pkg::*;
	import base_package::*;
	import obm_dut_cfg_package::*;
	`include "src/mac_tx_monitor.sv"
endpackage
import mac_tx_package::*;
