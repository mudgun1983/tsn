//PHY_PORT_TABLE
`define PHY_PORT_TABLE_STATUS	'h0020		
`define PHY_PORT_TABLE_CONTROL	'h0022	
`define PHY_PORT_TABLE_DIN_0	'h0024	
`define PHY_PORT_TABLE_DIN_1	'h0026
`define PHY_PORT_TABLE_DIN_2	'h0028
`define PHY_PORT_TABLE_DIN_3	'h002A
`define PHY_PORT_TABLE_DIN_4	'h002C
`define PHY_PORT_TABLE_DIN_5	'h002E
`define PHY_PORT_TABLE_DIN_6	'h0030

//LOGIC_PORT_TABLE	
`define LOGIC_PORT_TABLE_STATUS	 'h0200	
`define LOGIC_PORT_TABLE_CONTROL 'h0202	
`define LOGIC_PORT_TABLE_DIN_0	 'h0204	
`define LOGIC_PORT_TABLE_DIN_1	 'h0206
`define LOGIC_PORT_TABLE_DIN_2	 'h0208
`define LOGIC_PORT_TABLE_DIN_3	 'h020A
`define LOGIC_PORT_TABLE_DIN_4	 'h020C
`define LOGIC_PORT_TABLE_DIN_5	 'h020E
`define LOGIC_PORT_TABLE_DIN_6	 'h0210
`define LOGIC_PORT_TABLE_DIN_7	 'h0212
