library verilog;
use verilog.vl_types.all;
entity mac_pkg is
end mac_pkg;
