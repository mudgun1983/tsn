library verilog;
use verilog.vl_types.all;
entity pcs_env_pkg is
end pcs_env_pkg;
