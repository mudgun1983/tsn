library verilog;
use verilog.vl_types.all;
entity gmii_rx_if is
end gmii_rx_if;
