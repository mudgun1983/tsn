library verilog;
use verilog.vl_types.all;
entity xgmii64_tx_if is
end xgmii64_tx_if;
